`timescale 1ns / 1ps
`ifndef ONE // 1
`define ONE(WL) {{(WL-1){1'b0}}, 1'b1}
`endif

`ifndef ZERO // 0
`define ZERO(WL) {(WL){1'b0}}
`endif

`ifndef ALL1 // 111111
`define ALL1(WL) {(WL){1'b1}}
`endif

module Pipline_tb();

    parameter DATA_WL = 32'd32;
    parameter ADDR_WL = 32'd32;
    parameter WEA_WL  = 32'd4;
    parameter SW_ENV_NUM = 30'd320;
    parameter RAM_ADDR_WL = 12; // if RAM_ADDR_WL is 32, simulation will be very slow 

    reg        clk = 0;
    reg        rstn;
    reg [63:0] clk_cnt;
    reg [63:0] cycle_cnt;

    reg new_round; // a new round of compute is started

    // Pipeline ports
        wire [DATA_WL-1:0] uut_i_data;
        wire [DATA_WL-1:0] uut_o_data;
        wire [ADDR_WL-1:0] uut_o_addr;
        wire               uut_o_en;
        wire [WEA_WL-1:0]  uut_o_wea;
        wire               uut_o_rstb;

    // BRAM ports
        reg                    ram_i_wr1;
        reg  [RAM_ADDR_WL-1:0] ram_i_addr1;
        reg  [DATA_WL-1:0]     ram_i_data1;
        wire [DATA_WL-1:0]     ram_o_data1;
        wire                   ram_i_wr2;
        wire [RAM_ADDR_WL-1:0] ram_i_addr2;
        wire [DATA_WL-1:0]     ram_i_data2;
        wire [DATA_WL-1:0]     ram_o_data2;

    always #5 clk = !clk;

    initial begin
        rstn = 1;
        #10 rstn = 0;
        #10 rstn = 1;
    //  #10000 $finish;
    end

    always @(posedge clk or negedge rstn) begin
        if (rstn == 1'b0) begin
            clk_cnt <= 64'b0;
        end else begin
            clk_cnt <= clk_cnt + 1'b1;
        end
    end
    initial begin // write initial data
        #0  ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0; ram_i_data1 = 32'd0; new_round = 1'b0;
        // 1st round:
            #20 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'hb98e5284; // x0:-0.00027145829517394304
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'hbbf2b25e; // ẋ0:-0.007406516931951046
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h3d239cf2; // θ0:0.0399445965886116
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'hbbd215eb; // ω0:-0.006411304231733084

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'hbbc98439; // x1:-0.00614979537203908
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h3c1f3084; // ẋ1:0.009716156870126724
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'hbbe5d4bc; // θ1:-0.0070138853043317795
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'hbc484533; // ω1:-0.012223529629409313

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h3d428df8; // x2:0.0474986732006073
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'hbd23c960; // ẋ2:-0.03998696804046631
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'hbc3ec244; // θ2:-0.011642996221780777
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'hbc6168c4; // ω2:-0.013757888227701187

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h3bd45956; // x3:0.006480376236140728
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h3c4be384; // ẋ3:0.012444380670785904
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h3c8f7f0c; // θ3:0.017516635358333588
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'hb8c56a94; // ω3:-9.4135437393561e-05

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'hbccd9bbb; // x4:-0.02509867213666439
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'hbd38b506; // ẋ4:-0.04509451240301132
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h3cd2f202; // θ4:0.025750163942575455
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h3c9c758b; // ω4:0.01909901760518551

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h3d11388b; // x5:0.035454314202070236
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'hbd40dd6e; // ẋ5:-0.04708617180585861
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'hbd24498e; // θ5:-0.04010920971632004
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'hbd354503; // ω5:-0.04425526782870293

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'hbd2d0485; // x6:-0.04224063828587532
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'hbd485521; // ẋ6:-0.04890931025147438
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h3bda0097; // θ6:0.0066529023461043835
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h3d35e41a; // ω6:0.044406987726688385

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'hbba01cde; // x7:-0.004886253736913204
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'hbd2a658b; // ẋ7:-0.04160074517130852
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'hbb405969; // θ7:-0.0029350167606025934
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h3c8bc7f5; // ω7:0.017063120380043983

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h3d05d23a; // x8:0.03267119079828262
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h3cfcd970; // ẋ8:0.030865401029586792
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'hba9ec12f; // θ8:-0.001211201655678451
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'hbc2c89c0; // ω8:-0.01053088903427124

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h3c99b1b5; // x9:0.018761495128273964
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'hbd45630a; // ẋ9:-0.0481901541352272
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h3c39a724; // θ9:0.011331353336572647
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'hbcd631e9; // ω9:-0.026146845892071724

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h3c3fb4ce; // x10:0.011700822040438652
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'hbbd73515; // ẋ10:-0.006567607168108225
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h3d012767; // θ10:0.031531717628240585
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'hb9c72450; // ω10:-0.0003798329271376133

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'hbc1bfbb1; // x11:-0.009520457126200199
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h3c0f3437; // ẋ11:0.008740476332604885
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'hbcc85f08; // θ11:-0.02445937693119049
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h3cc4a8be; // ω11:0.02400624379515648

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h3c5eba32; // x12:0.013594197109341621
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h3c3b7e17; // ẋ12:0.011443636380136013
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h3d36dfa1; // θ12:0.044646862894296646
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'hbc79296c; // ω12:-0.015207629650831223

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'hbcb1df72; // x13:-0.02171299234032631
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'hbcf5a2a6; // ẋ13:-0.02998478338122368
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h3d30ad96; // θ13:0.04313429445028305
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'hbc6eaef6; // ω13:-0.014568081125617027

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'hbcd27152; // x14:-0.02568880096077919
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h3d40efec; // ẋ14:0.04710380733013153
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h3d2468da; // θ14:0.040139056742191315
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'hbd263817; // ω14:-0.040580835193395615

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'hbd0a47e3; // x15:-0.033759962767362595
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h3c41c806; // ẋ15:0.01182747446000576
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h3bfc2cef; // θ15:0.007695786189287901
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'hbc149f91; // ω15:-0.009071246720850468

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h3adcf5c7; // x16:0.001685791532509029
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h3cb15c2c; // ẋ16:0.021650396287441254
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'hbc28061f; // θ16:-0.010255365632474422
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h3cec8795; // ω16:0.028873244300484657

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h3bf18013; // x17:0.007370003964751959
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h3a5f657c; // ẋ17:0.0008521897252649069
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'hbb03f5e6; // θ17:-0.002013558056205511
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h3d0b1aca; // ω17:0.03396109491586685

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'hbc884336; // x18:-0.016633611172437668
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h3ce29752; // ẋ18:0.02766004577279091
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h3d0307ad; // θ18:0.03198974207043648
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'hbc1ee223; // ω18:-0.009697469882667065

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h3cc27bde; // x19:0.023740705102682114
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h3cfc3cc0; // ẋ19:0.03079068660736084
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'hbca6787c; // θ19:-0.02032112330198288
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'hbcf0fe27; // ω19:-0.029418064281344414

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'hbd2b0732; // x20:-0.04175490885972977
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h3c9edac8; // ẋ20:0.019391432404518127
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'hbc0ea232; // θ20:-0.008705662563443184
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h3c0c6a57; // ω20:0.008570275269448757

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h3c075497; // x21:0.008259913884103298
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h3cd77883; // ẋ21:0.026302581652998924
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h3bcd9a8c; // θ21:0.006274526938796043
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'hb967198f; // ω21:-0.00022039398027118295

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h3c37729c; // x22:0.011196758598089218
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'hbd2e66c1; // ẋ22:-0.04257846251130104
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'hbc54f05f; // θ22:-0.012996762059628963
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h3c7c0cf9; // ω22:0.015383952297270298

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h3bc550db; // x23:0.006021601613610983
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'hbb89e523; // ẋ23:-0.004208223428577185
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h3d233866; // θ23:0.03984870761632919
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h3ca9a3bd; // ω23:0.020707959309220314

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'hb920c531; // x24:-0.0001533224858576432
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'hbd28af9d; // ẋ24:-0.04118310287594795
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'hbcfa6645; // θ24:-0.030566344037652016
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h3d25f9a4; // ω24:0.040521278977394104

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'hbd1a620c; // x25:-0.037691161036491394
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'hbc484852; // ẋ25:-0.012224273756146431
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'hbad10434; // θ25:-0.0015946687199175358
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h396b9d98; // ω25:0.00022470054682344198

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h3ce87120; // x26:0.02837425470352173
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'hbd15b196; // ẋ26:-0.036546312272548676
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h3c5944e3; // θ26:0.013261052779853344
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h3be69259; // ω26:0.0070364889688789845

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'hbcb537cb; // x27:-0.022121330723166466
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h3d3de56a; // ẋ27:0.04636136442422867
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h3a97f9c9; // θ27:0.0011594827519729733
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'hbd395f87; // ω27:-0.045257117599248886

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h3c444c73; // x28:0.0119811175391078
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h3c1d67d9; // ẋ28:0.009607278741896152
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'hbd1764e9; // θ28:-0.03696146979928017
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'hbcf989de; // ω28:-0.030461248010396957

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h3bb92e2a; // x29:0.005651255138218403
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h3c24c31b; // ẋ29:0.01005628239363432
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h3d1b57e8; // θ29:0.03792563080787659
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h3d43bba6; // ω29:0.04778637737035751

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h3c215a44; // x30:0.009848181158304214
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'hbc92c341; // ẋ30:-0.01791536994278431
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'hbcda6385; // θ30:-0.026658782735466957
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h3c61ffb1; // ω30:0.013793871738016605

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h3b16ed55; // x31:0.002302964450791478
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h3c89c1e6; // ẋ31:0.016816090792417526
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h3d187d04; // θ31:0.037228599190711975
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h3b92cb68; // ω31:0.004479814320802689

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h3ca7cc56; // x32:0.02048317715525627
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'hbcf9ae05; // ẋ32:-0.03047848679125309
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h3ced1e40; // θ32:0.028945088386535645
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h3c6cd1f3; // ω32:0.014454352669417858

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h3d38adc8; // x33:0.045087605714797974
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h3d1491e6; // ẋ33:0.03627195209264755
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'hbce0c2f8; // θ33:-0.027436718344688416
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h3d1e6131; // ω33:0.03866690769791603

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h3c4c8905; // x34:0.012483839876949787
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'hbcb539dc; // ẋ34:-0.02212231606245041
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h3d16bfc1; // θ34:0.0368039645254612
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'hbc96d625; // ω34:-0.01841265894472599

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h3d28cfe5; // x35:0.04121388867497444
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'hbcb06614; // ẋ35:-0.021533049643039703
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'hbd32ac2e; // θ35:-0.043621234595775604
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h3c3c4c24; // ω35:0.011492762714624405

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'hbcae9827; // x36:-0.021312786266207695
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h3a464e0c; // ẋ36:0.0007564730476588011
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'hbc2d522d; // θ36:-0.010578674264252186
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h3ca06469; // ω36:0.019579129293560982

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'hb953630d; // x37:-0.00020159427367616445
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h3cafdf9c; // ẋ37:0.021468929946422577
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h3bf5543e; // θ37:0.007486849091947079
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h3d35779f; // ω37:0.0443035326898098

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h3d29de7a; // x38:0.0414719358086586
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h3cb04d84; // ẋ38:0.02152133733034134
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h3ce6ab13; // θ38:0.02815774641931057
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h3d4a3ca2; // ω38:0.049374230206012726

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'hbd182c54; // x39:-0.037151649594306946
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h3d2c0816; // ẋ39:0.041999898850917816
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'hbc079ebe; // θ39:-0.008277593180537224
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'hbcfa6c5d; // ω39:-0.030569249764084816

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'hbbaacf0e; // x40:-0.005212671123445034
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h3d06a7bc; // ẋ40:0.032874807715415955
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'hbc97c82a; // θ40:-0.018528062850236893
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'hbd3c2b07; // ω40:-0.04593947157263756

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'hbc59073e; // x41:-0.013246355578303337
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'hbab935c9; // ẋ41:-0.001413040910847485
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'hbcabe9cb; // θ41:-0.020985504612326622
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'hbce25596; // ω41:-0.02762870118021965

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'hbcbdad9f; // x42:-0.02315407805144787
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h3cdb05cf; // ẋ42:0.026736168190836906
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h3a81fd31; // θ42:0.0009917375864461064
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h3ca5ae6d; // ω42:0.02022477425634861

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h3ca90961; // x43:0.020634355023503304
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'hbbb608cb; // ẋ43:-0.00555524742230773
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'hbbd98a21; // θ43:-0.006638780701905489
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'hbd32a94e; // ω43:-0.043618492782115936

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'hbd1a2a90; // x44:-0.03763824701309204
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'hbc47fbcd; // ẋ44:-0.012206030078232288
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h3cd31844; // θ44:0.025768406689167023
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h3c82a2d1; // ω44:0.015946777537465096

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'hbcc02522; // x45:-0.02345520630478859
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'hbb732805; // ẋ45:-0.003710271092131734
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h3c8f04d8; // θ45:0.017458364367485046
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h3d0e03ec; // ω45:0.034671708941459656

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h3d4365a6; // x46:0.047704361379146576
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'hbc622f1f; // ẋ46:-0.013805179856717587
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'hbd36ec74; // θ46:-0.0446590930223465
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h3c90e0d5; // ω46:0.017685333266854286

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'hbc9fcb30; // x47:-0.019506067037582397
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'hbce05fe3; // ẋ47:-0.027389472350478172
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'hbcdcf5c0; // θ47:-0.026972651481628418
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h3c71084c; // ω47:0.014711450785398483

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h3ca1570e; // x48:0.01969483122229576
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'hbc9f5814; // ẋ48:-0.01945117861032486
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h3d3baa13; // θ48:0.04581649228930473
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h3d02ba15; // ω48:0.03191574290394783

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h3c7ad39b; // x49:0.015309239737689495
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h3c4b1ea0; // ẋ49:0.012397438287734985
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h3b50881f; // θ49:0.0031819415744394064
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'hbca28181; // ω49:-0.019837142899632454

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'hbcca3bc5; // x50:-0.024686703458428383
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'hbd1adac3; // ẋ50:-0.03780628368258476
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'hbcf40a86; // θ50:-0.029790174216032028
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'hba0396a1; // ω50:-0.0005019698874093592

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h3cd919a7; // x51:0.026501489803195
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h3c208535; // ẋ51:0.009797384031116962
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'hbc72b554; // θ51:-0.01481373980641365
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'hbc6d0798; // ω51:-0.014467142522335052

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'hbc809d02; // x52:-0.01569986715912819
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'hbc6f2277; // ẋ52:-0.014595619402825832
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h3cfe85cf; // θ52:0.031069664284586906
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'hbcd42263; // ω52:-0.02589530311524868

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'hbb95547d; // x53:-0.004557190928608179
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h3d47496b; // ẋ53:0.04865400120615959
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'hbbe314fc; // θ53:-0.006929991766810417
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'hbc8645e5; // ω53:-0.01639075018465519

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'hbc0bb491; // x54:-0.0085269371047616
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h3d49f50a; // ẋ54:0.049305953085422516
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'hb95c33a2; // θ54:-0.00021000069682486355
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'hbd27dd3e; // ω54:-0.040982477366924286

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'hbcf97b7e; // x55:-0.030454393476247787
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h3cef83b1; // ẋ55:0.029237600043416023
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'hbd032ac4; // θ55:-0.03202320635318756
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h3bb13c15; // ω55:0.00540877366438508

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h3cf9b9d8; // x56:0.030484125018119812
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'hbd053e48; // ẋ56:-0.03253009915351868
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'hbcb4e59a; // θ56:-0.022082138806581497
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h3ce633ee; // ω56:0.028100933879613876

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h3c57f8f1; // x57:0.01318191085010767
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h3d37b47a; // ẋ57:0.04484985023736954
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h3ca20d53; // θ57:0.019781744107604027
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h3d46dff0; // ω57:0.048553407192230225

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h3d363b6d; // x58:0.0444902665913105
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h3c836a12; // ẋ58:0.016041789203882217
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h3b2c537c; // θ58:0.0026294877752661705
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h3d0dcd0c; // ω58:0.03461937606334686

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'hbd073334; // x59:-0.03300781548023224
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h3c9e6127; // ẋ59:0.019333435222506523
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'hbcc1a150; // θ59:-0.02363649010658264
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'hbd2209c7; // ω59:-0.03956010565161705

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'hbbda66db; // x60:-0.0066650933586061
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h3b0331ab; // ẋ60:0.002001861808821559
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'hbaf9416f; // θ60:-0.001901669311337173
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'hbb63870d; // ω60:-0.0034717947710305452

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h3d1e4edf; // x61:0.038649436086416245
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'hbba479d2; // ẋ61:-0.005019404925405979
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h3ca1b0c6; // θ61:0.019737612456083298
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'hbb94b35b; // ω61:-0.004537982400506735

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h3bd2c3c1; // x62:0.006432027090340853
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h3ab04b26; // ẋ62:0.0013450130354613066
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'hbc6b7d7d; // θ62:-0.014373180456459522
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h3b76a116; // ω62:0.0037632635794579983

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'hbcc889ee; // x63:-0.024479832500219345
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h3d36bb9a; // ẋ63:0.04461250454187393
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'hbd0034d7; // θ63:-0.031300392001867294
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'hbcf64ad2; // ω63:-0.03006497398018837

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'hbc91cd66; // x64:-0.017798136919736862
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h3bc08aa9; // ẋ64:0.005875904578715563
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'hbaa0d095; // θ64:-0.0012269193539395928
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'hbc80a229; // ω64:-0.015702323988080025

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h3c4b6f86; // x65:0.012416725978255272
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h3d13c7d1; // ẋ65:0.03607923164963722
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h3c46030d; // θ65:0.012085688300430775
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'hbc8fdf70; // ω65:-0.01756259799003601

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h3c7d5ee8; // x66:0.015464521944522858
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'hbc28a283; // ẋ66:-0.010292652063071728
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h3d202c31; // θ66:0.0391046442091465
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'hbc20c4ea; // ω66:-0.009812572970986366

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'hbd0b7c84; // x67:-0.03405429422855377
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h3bd2f08a; // ẋ67:0.006437365896999836
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'hbc576cb7; // θ67:-0.013148478232324123
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h3beb0893; // ω67:0.0071726529859006405

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h3d19792d; // x68:0.03746907785534859
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h39d5e965; // ẋ68:0.0004080041835550219
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'hbc4da084; // θ68:-0.0125504769384861
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'hbd42ab83; // ω68:-0.04752684757113457

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h3d17f835; // x69:0.03710194304585457
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h3c81b24b; // ẋ69:0.01583208702504635
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h3cc591b5; // θ69:0.024117330089211464
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h3c4e18a3; // ω69:0.0125791160389781

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h3d29031e; // x70:0.04126273840665817
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h3d108c4b; // ẋ70:0.03529004380106926
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h3d41b393; // θ70:0.04729039594531059
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h3d2a757d; // ω70:0.04161595180630684

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h3cec0520; // x71:0.02881103754043579
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h3d248e69; // ẋ71:0.040174875408411026
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'hbd35b2da; // θ71:-0.04436001926660538
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h3c7160e9; // ω71:0.014732577838003635

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'hbca17970; // x72:-0.019711226224899292
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'hbc4b29e1; // ẋ72:-0.012400121428072453
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h3cce53b0; // θ72:0.025186389684677124
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'hbb72cbd5; // ω72:-0.0037047762889415026

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'hbccd0d3b; // x73:-0.025030722841620445
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'hbc843ad1; // ẋ73:-0.01614132709801197
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h3c9d3223; // θ73:0.01918894611299038
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h3cee5597; // ω73:0.0290935467928648

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h3cb570b2; // x74:0.022148463875055313
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h3c0b4d3b; // ẋ74:0.008502299897372723
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h3c3a8d5e; // θ74:0.011386243626475334
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h3cdf34da; // ω74:0.027246881276369095

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'hbc8d9e1d; // x75:-0.01728730835020542
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h3cd524aa; // ẋ75:0.026018459349870682
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h3d00c21d; // θ75:0.03143512085080147
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'hbc486653; // ω75:-0.012231427244842052

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h3d18e354; // x76:0.03732617199420929
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h3d4b1e2f; // ẋ76:0.049589332193136215
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h3ce36db7; // θ76:0.02776227705180645
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'hbd47c0a6; // ω76:-0.048767708241939545

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h3c28720b; // x77:0.010281096212565899
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h3d3f9521; // ẋ77:0.04677307978272438
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h3d3bf048; // θ77:0.04588344693183899
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'hbb3634a0; // ω77:-0.002780236303806305

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'hbcee77b4; // x78:-0.029109813272953033
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h3d0a10f0; // ẋ78:0.03370755910873413
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h3d25adfa; // θ78:0.0404491201043129
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'hbb89df1c; // ω78:-0.004207504913210869

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h3d14a806; // x79:0.03629305213689804
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h3caba8ed; // ẋ79:0.020954573526978493
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'hbd1b99bf; // θ79:-0.03798842057585716
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'hbd37a53a; // ω79:-0.04483530670404434

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h3ca49dc9; // x80:0.020094769075512886
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h3c0ced75; // ẋ80:0.0086015360429883
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h3c08d8d0; // θ80:0.008352473378181458
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'hbc59124e; // ω80:-0.013248993083834648

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'hbca0d459; // x81:-0.019632505252957344
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h3b5d4100; // ẋ81:0.0033760666847229004
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'hbcbb1020; // θ81:-0.022834837436676025
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'hbc204d7c; // ω81:-0.009784098714590073

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'hbd0c821b; // x82:-0.03430376574397087
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'hbc7905d9; // ẋ82:-0.0151991480961442
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'hba90b711; // θ82:-0.0011040886165574193
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'hbc8139a7; // ω82:-0.0157745610922575

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h3c70c92b; // x83:0.014696399681270123
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'hbc1c6a3a; // ẋ83:-0.009546810761094093
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h3ce5d1e2; // θ83:0.02805418148636818
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'hbc633306; // ω83:-0.013867145404219627

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'hbd42279b; // x84:-0.047401051968336105
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h3ceb5d9a; // ẋ84:0.028731156140565872
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h39fa2690; // θ84:0.0004771244712173939
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'hbd32a61e; // ω84:-0.04361545294523239

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'hbd3e2614; // x85:-0.04642303287982941
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h3d2ec03c; // ẋ85:0.04266379773616791
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'hbd201886; // θ85:-0.039085887372493744
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h3cf2dfd5; // ω85:0.029647747054696083

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'hbd3d86fb; // x86:-0.04627130553126335
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'hbcbebd6a; // ẋ86:-0.02328367903828621
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'hbc6e772d; // θ86:-0.014554780907928944
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h3cbd8361; // ω86:0.023133935406804085

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h3cf95fad; // x87:0.030441129580140114
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'hbd25de88; // ẋ87:-0.04049542546272278
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'hbd0b2356; // θ87:-0.033969245851039886
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'hbd28464b; // ω87:-0.04108266159892082

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'hbc9821dc; // x88:-0.018570832908153534
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h3cb8c062; // ẋ88:0.022552672773599625
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h3caa4696; // θ88:0.020785611122846603
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h3d48bce6; // ω88:0.04900827258825302

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h3c936283; // x89:0.017991309985518456
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h3cb45cb3; // ẋ89:0.0220168586820364
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'hbc3bca04; // θ89:-0.011461738497018814
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h3d222da8; // ω89:0.03959432244300842

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h3d29ee5a; // x90:0.04148707538843155
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h3bd886ff; // ẋ90:0.006607889663428068
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h3d42848d; // θ90:0.04748969152569771
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h3b447c5f; // ω90:0.0029981357511132956

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h3d10f7a3; // x91:0.03539241477847099
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'hbce31879; // ẋ91:-0.027721630409359932
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h3cb73849; // θ91:0.02236570604145527
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'hbd03acb6; // ω91:-0.032147131860256195

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'hbd107d49; // x92:-0.03527573123574257
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'hbcf41dcd; // ẋ92:-0.029799366369843483
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h3d1a5ccd; // θ92:0.03768615797162056
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'hbc89b9c5; // ω92:-0.016812214627861977

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h3ce5efbc; // x93:0.028068415820598602
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'hbd21f125; // ẋ93:-0.03953661397099495
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'hbcfac7a3; // θ93:-0.030612772330641747
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h3cee3bc2; // ω93:0.029081229120492935

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h3c6d932b; // x94:0.014500419609248638
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'hbcfc2ebe; // ẋ94:-0.030784007161855698
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h3c23af6a; // θ94:0.009990552440285683
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'hbad60730; // ω94:-0.0016329046338796616

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h3d27b43b; // x95:0.040943365544080734
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'hbbc70f2e; // ẋ95:-0.006074807606637478
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h3d195df8; // θ95:0.0374431312084198
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h3d29716d; // ω95:0.04136793687939644

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h3d37077a; // x96:0.044684864580631256
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'hbb090e68; // ẋ96:-0.0020913127809762955
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3a8bfe25; // θ96:0.0010680599370971322
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3d324c4b; // ω96:0.04352978989481926

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3d319a50; // x97:0.04336005449295044
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbb162c3e; // ẋ97:-0.0022914553992450237
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3c7f5cc2; // θ97:0.01558608002960682
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbce4ce2a; // ω97:-0.02793033793568611

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'hbce72aea; // x98:-0.02821870520710945
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h3cfc3725; // ẋ98:0.030788013711571693
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'hbc71ecb4; // θ98:-0.0147659070789814
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbd43282b; // ω98:-0.047645729035139084

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'hbcd741bb; // x99:-0.02627645991742611
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbd49b2fd; // ẋ99:-0.04924296215176582
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h3ce640f2; // θ99:0.028107140213251114
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3c81b791; // ω99:0.01583460159599781

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'hbcef7455; // x100:-0.029230276122689247
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h3d3f692b; // ẋ100:0.04673115536570549
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'hbcd8be9b; // θ100:-0.026458075270056725
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbd2821fc; // ω100:-0.04104803502559662

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'hbcb0d31e; // x101:-0.021585043519735336
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbd3bafd5; // ẋ101:-0.045821983367204666
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'hbcd6a371; // θ101:-0.026200981810688972
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbca6a1fe; // ω101:-0.020340915769338608

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h3d24bcd3; // x102:0.04021913930773735
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3d010437; // ẋ102:0.03149816021323204
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h3ccf0709; // θ102:0.025271909311413765
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'hbc0d2615; // ω102:-0.008615036495029926

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'hbd080f3a; // x103:-0.033217646181583405
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h3c81b0e9; // ẋ103:0.01583142764866352
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3d068a86; // θ103:0.032846949994564056
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbb9dee26; // ω103:-0.004819649271667004

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbc859ad4; // x104:-0.016309179365634918
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3d0c34f5; // ẋ104:0.03423019126057625
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h3d1f535b; // θ104:0.03889785334467888
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3d03b446; // ω104:0.03215434402227402

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3d390338; // x105:0.04516908526420593
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h3c63844d; // ẋ105:0.013886523433029652
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbc826730; // θ105:-0.015918344259262085
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'hbd14869d; // ω105:-0.036261189728975296

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3ca3dcd0; // x106:0.020002752542495728
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbc984d31; // ẋ106:-0.018591495230793953
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'hbd10fb79; // θ106:-0.03539607301354408
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbb354e2f; // ω106:-0.002766500925645232

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3d1ddea0; // x107:0.03854238986968994
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'hbc9f7b71; // ẋ107:-0.019468041136860847
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbb247a1f; // θ107:-0.002509720390662551
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'hbcaa8518; // ω107:-0.020815417170524597

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'hbcf4dd6a; // x108:-0.02989073470234871
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbce8721f; // ẋ108:-0.028374729678034782
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbc00ac88; // θ108:-0.007853634655475616
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbc182da7; // ω108:-0.009288228116929531

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h3c8f1c63; // x109:0.01746959052979946
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h3cdb32ca; // ẋ109:0.0267576165497303
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'hbc59635b; // θ109:-0.013268317095935345
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h3caab71c; // ω109:0.02083926647901535

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h3d0e341e; // x110:0.03471767157316208
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbd045242; // ẋ110:-0.03230500966310501
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3cc294a2; // θ110:0.023752514272928238
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'hbc5bb06e; // ω110:-0.013408763334155083

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbd3d8eff; // x111:-0.046278949826955795
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3cea98c1; // ẋ111:0.028637291863560677
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3d379e98; // θ111:0.044828981161117554
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'hbd386ecf; // ω111:-0.04502755030989647

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'hbd25fe99; // x112:-0.04052600637078285
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3b5f6bec; // ẋ112:0.003409142605960369
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbaa23501; // θ112:-0.0012375415535643697
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbc267b48; // ω112:-0.010161228477954865

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'hbd475050; // x113:-0.04866057634353638
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3d457702; // ẋ113:0.04820919781923294
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h3c5eda88; // θ113:0.013601906597614288
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'hbc150681; // ω113:-0.009095788933336735

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'hbba6786b; // x114:-0.005080272909253836
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3d167ff5; // ẋ114:0.03674312308430672
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3ce239f5; // θ114:0.02761552669107914
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'hbcb25a40; // ω114:-0.021771550178527832

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'hbc72d883; // x115:-0.014822128228843212
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h3d0265a0; // ẋ115:0.031835198402404785
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbcb0edf7; // θ115:-0.021597845479846
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbd3356fd; // ω115:-0.04378413036465645

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3cc71a09; // x116:0.024304406717419624
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'hbc06d35c; // ẋ116:-0.008229102939367294
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h3d362f94; // θ116:0.044478967785835266
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h3cc35456; // ω116:0.023843925446271896

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbc5382b2; // x117:-0.012909578159451485
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbcbddfdd; // ẋ117:-0.023178035393357277
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'hbcd5e2a6; // θ117:-0.02610905095934868
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'hbd0b127e; // ω117:-0.03395318239927292

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbd07f2fa; // x118:-0.03319070488214493
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h3c34a80e; // ẋ118:0.011026395484805107
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'hbcac2f58; // θ118:-0.02101866900920868
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3cdd802d; // ω118:0.027038658037781715

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h3d022643; // x119:0.031774770468473434
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h3d3b4945; // ẋ119:0.04572417214512825
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'hbc860906; // θ119:-0.016361724585294724
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h3d1c6165; // ω119:0.03817882016301155

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h3cd5a660; // x120:0.026080310344696045
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'hbccca007; // ẋ120:-0.024978650733828545
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h3d4208eb; // θ120:0.04737178608775139
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'hbcca57bc; // ω120:-0.024700038135051727

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'hbd1b3f76; // x121:-0.03790231794118881
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h3d05365f; // ẋ121:0.03252255544066429
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3b6d95c7; // θ121:0.0036252604331821203
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbb712f8b; // ω121:-0.0036802019458264112

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'hbc913f23; // x122:-0.01773030124604702
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h3d24f62c; // ẋ122:0.04027383029460907
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3d3f132c; // θ122:0.04664914309978485
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbd1c517c; // ω122:-0.038163647055625916

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3cde5956; // x123:0.027142208069562912
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'hbc936ffd; // ẋ123:-0.017997736111283302
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h3cccf0db; // θ123:0.02501719258725643
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h3ce35095; // ω123:0.027748385444283485

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3c328e26; // x124:0.010898148640990257
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h3c01ca65; // ẋ124:0.007921789772808552
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h3cefb67c; // θ124:0.029261820018291473
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'hbca5b6c2; // ω124:-0.02022874727845192

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'hbca54b21; // x125:-0.02017742581665516
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3ca936b4; // ẋ125:0.02065596729516983
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'hbd1e173c; // θ125:-0.03859637677669525
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3cb30960; // ω125:0.021855056285858154

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h3d0f5c68; // x126:0.035000234842300415
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3c93cf4c; // ẋ126:0.01804318279027939
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h3d123206; // θ126:0.0356922373175621
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3cd7297c; // ω126:0.026264898478984833

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3c25d37d; // x127:0.010121223516762257
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h3d1fb4a3; // ẋ127:0.038990627974271774
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbcd0e50a; // θ127:-0.025499839335680008
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3bdbc0ab; // ω127:0.00670631742104888

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h3cb30daa; // x128:0.02185710147023201
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'hbc7985a4; // ẋ128:-0.015229616314172745
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'hbc3bf86d; // θ128:-0.01147280354052782
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbd1562ce; // ω128:-0.036471180617809296

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h3d4a04dd; // x129:0.049321044236421585
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3cf857ce; // ẋ129:0.030315306037664413
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3aa6a3c6; // θ129:0.001271360320970416
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'hbbf9c6bc; // ω129:-0.0076225679367780685

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'hbd46ead1; // x130:-0.04856378212571144
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'hbc0a4321; // ẋ130:-0.008438856340944767
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'hbcb7b9b8; // θ130:-0.022427424788475037
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'hbc8355ee; // ω130:-0.016032185405492783

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'hbc1f3667; // x131:-0.00971756037324667
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h3c801540; // ẋ131:0.015635132789611816
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'hbd1c9b8f; // θ131:-0.03823428973555565
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h3c8f98dd; // ω131:0.017528945580124855

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3caeac42; // x132:0.021322373300790787
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'hbc01e65b; // ẋ132:-0.00792845617979765
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'hbd3e7fcf; // θ132:-0.046508606523275375
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbcc47fcf; // ω132:-0.023986725136637688

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'hbc915b1f; // x133:-0.01774364523589611
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h3d3e5095; // ẋ133:0.04646356776356697
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'hbcb706b3; // θ133:-0.02234206162393093
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbcbbbd6b; // ω133:-0.02291746996343136

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'hbc8e8fe8; // x134:-0.01740260422229767
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3cbff972; // ẋ134:0.02343437448143959
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h3c88fb02; // θ134:0.016721252351999283
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h3d4be458; // ω134:0.04977831244468689

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h3d469cbf; // x135:0.04848932847380638
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbbd1327e; // ẋ135:-0.00638419296592474
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h3d0d5c03; // θ135:0.03451157733798027
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h3d38ae4b; // ω135:0.04508809372782707

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbcb55309; // x136:-0.022134320810437202
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'hbc69d579; // ẋ136:-0.014272087253630161
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'hbc03ee70; // θ136:-0.008052453398704529
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h3cee6a74; // ω136:0.029103495180606842

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h3d21393d; // x137:0.03936122730374336
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'hbd172fa0; // ẋ137:-0.03691065311431885
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h3b9745fa; // θ137:0.004616496153175831
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbc4379ad; // ω137:-0.011930865235626698

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3d0623b0; // x138:0.03274887800216675
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbbcb872b; // ẋ138:-0.00621118163689971
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h3cdcdca0; // θ138:0.026960670948028564
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'hbd36e910; // ω138:-0.04465585947036743

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3a784ea5; // x139:0.0009472168167121708
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'hbd45d136; // ẋ139:-0.04829522222280502
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'hbd4a39da; // θ139:-0.04937157779932022
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3b5b9341; // ω139:0.00335045182146132

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'hbc22e844; // x140:-0.009943071752786636
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h3d21d073; // ẋ140:0.03950543329119682
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbc43b24b; // θ140:-0.011944363825023174
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h3c7aa3a9; // ω140:0.015297808684408665

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'hbcb7d3d5; // x141:-0.022439876571297646
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbc14d536; // ẋ141:-0.009084036573767662
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h3c0b7038; // θ141:0.008510641753673553
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h3c1d5c3b; // ω141:0.009604508988559246

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'hbd3e0d6f; // x142:-0.04639953002333641
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbc654d0c; // ẋ142:-0.013995420187711716
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3d1af489; // θ142:0.037830863147974014
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h3ce2d19d; // ω142:0.027687842026352882

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbd415b20; // x143:-0.04720604419708252
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbd4cc716; // ẋ143:-0.04999455064535141
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'hbcdbeb86; // θ143:-0.02684570476412773
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h3ae12ac2; // ω143:0.0017178880516439676

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'hbce486c1; // x144:-0.02789628691971302
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'hbd183e3f; // ẋ144:-0.03716873750090599
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'hbc06855c; // θ144:-0.008210506290197372
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h3bcc8b4b; // ω144:0.006242190953344107

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h3c35202c; // x145:0.011055033653974533
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h3d345363; // ẋ145:0.044024836272001266
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'hbd18d838; // θ145:-0.037315577268600464
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h3d195b61; // ω145:0.03744066134095192

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h3c17645b; // x146:0.009240235202014446
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'hbcfdbc65; // ẋ146:-0.03097362257540226
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'hbd06d5fa; // θ146:-0.03291890770196915
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h3c8f16b3; // ω146:0.01746687851846218

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'hbcfbbaf6; // x147:-0.030728798359632492
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h3ca6ef33; // ẋ147:0.020377730950713158
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'hbd2a3818; // θ147:-0.04155740141868591
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'hbd33da61; // ω147:-0.04390943422913551

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'hbd0ac1c6; // x148:-0.0338762030005455
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'hbb50b563; // ẋ148:-0.0031846396159380674
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h3d095386; // θ148:0.03352691978216171
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h3d001c41; // ω148:0.031276945024728775

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'hbcfe36fe; // x149:-0.031032081693410873
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'hbd379633; // ẋ149:-0.04482097551226616
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h3ccd03b1; // θ149:0.025026174262166023
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'hbc9d77d9; // ω149:-0.019222186878323555

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'hbb645ae5; // x150:-0.003484421642497182
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h3cbc2c06; // ẋ150:0.022970210760831833
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h3cb96da2; // θ150:0.022635284811258316
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'hbce4b08c; // ω150:-0.027916215360164642

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h3c897aef; // x151:0.016782252117991447
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'hbd44c9c2; // ẋ151:-0.04804397374391556
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'hbcac6739; // θ151:-0.021045314148068428
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'hbc9e29c8; // ω151:-0.019307032227516174

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h3d4c1732; // x152:0.04982680827379227
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'hbc9e2585; // ẋ152:-0.019305000081658363
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h3d23ad25; // θ152:0.039960045367479324
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'hbd071d71; // ω152:-0.03298706188797951

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'hbc001935; // x153:-0.007818509824573994
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h3d34360a; // ẋ153:0.04399684816598892
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'hbc603d1e; // θ153:-0.013686446473002434
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'hbca00ef7; // ω153:-0.019538385793566704

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'hbd0e353f; // x154:-0.034718748182058334
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h3cff2b52; // ẋ154:0.03114858642220497
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'hbd2bb82b; // θ154:-0.041923683136701584
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h3cd6b58d; // ω154:0.026209617033600807

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'hbc93b7e1; // x155:-0.01803201623260975
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'hbb131f04; // ẋ155:-0.0022448906674981117
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h3d395414; // θ155:0.045246198773384094
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h3c2f801c; // ω155:0.01071169599890709

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'hba9637e3; // x156:-0.001146074733696878
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'hbcbdf1ba; // ẋ156:-0.02318655326962471
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'hbd22ae88; // θ156:-0.03971722722053528
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h3b9bc835; // ω156:0.0047540911473333836

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'hbd26c5a7; // x157:-0.040715839713811874
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'hbd30ee81; // ẋ157:-0.04319620504975319
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'hbc7be41f; // θ157:-0.01537421252578497
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'hbb2f3b18; // ω157:-0.0026738103479146957

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'hbafbccb1; // x158:-0.0019210783066228032
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'hbb87ef9b; // ẋ158:-0.004148436244577169
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h3ca777ba; // θ158:0.02044283226132393
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h3c819c7f; // ω158:0.01582169346511364

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'hbd3e1428; // x159:-0.046405941247940063
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'hbd37d402; // ẋ159:-0.04487992078065872
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h3d1cb57c; // θ159:0.03825901448726654
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'hbd296c0a; // ω159:-0.04136279970407486

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h3d2acccc; // x160:0.04169921576976776
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h3d228bbb; // ẋ160:0.03968403860926628
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'hbc6df579; // θ160:-0.014523857273161411
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'hbd2de30c; // ω160:-0.0424528568983078

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h3b6d026c; // x161:0.0036164773628115654
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h3c8b403f; // ẋ161:0.0169984083622694
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'hbc0a95b8; // θ161:-0.008458547294139862
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h3cc4aad5; // ω161:0.024007240310311317

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h3ced5001; // x162:0.0289688128978014
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h3c9bced5; // ẋ162:0.01901952363550663
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h3ca2dfd0; // θ162:0.019882112741470337
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h3ce387b4; // ω162:0.027774669229984283

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h3d24d900; // x163:0.040246009826660156
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'hbd21fbf0; // ẋ163:-0.0395469069480896
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'hbd37252d; // θ163:-0.04471318796277046
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h3cb22d43; // ω163:0.02175009809434414

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'hbd121ca8; // x164:-0.03567185997962952
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'hbcf5e774; // ẋ164:-0.030017592012882233
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h3d39513d; // θ164:0.04524349048733711
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'hbcd3a3b4; // ω164:-0.02583489567041397

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'hbcad20a2; // x165:-0.021133724600076675
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h3d2288f6; // ẋ165:0.03968139737844467
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h3ae743b1; // θ165:0.001764407497830689
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'hbcda52e4; // ω165:-0.02665085345506668

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'hbc37f06e; // x166:-0.011226756498217583
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h3b4aea7e; // ẋ166:0.003096252214163542
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'hbb92fe2c; // θ166:-0.00448586605489254
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h3cde2313; // ω166:0.027116334065794945

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h3d066c2c; // x167:0.03281800448894501
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h3b9ddcc7; // ẋ167:0.004817578475922346
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h3cc5f12b; // θ167:0.02416284941136837
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'hba8efcdb; // ω167:-0.0010909097036346793

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h3ab469bc; // x168:0.0013764421455562115
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h3d42d37d; // ẋ168:0.047564972192049026
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h3c0faa91; // θ168:0.008768693543970585
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h3cf8641e; // ω168:0.03032117709517479

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'hbc79c39c; // x169:-0.015244390815496445
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'hbd21512a; // ẋ169:-0.03938404470682144
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h3c83e5d3; // θ169:0.016100799664855003
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h3c61fe67; // ω169:0.013793564401566982

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'hbd332185; // x170:-0.0437331385910511
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h3caf1aab; // ẋ170:0.0213750209659338
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'hbc520903; // θ170:-0.012819531373679638
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h3ca4b677; // ω170:0.020106537267565727

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h3d28f4c7; // x171:0.04124906286597252
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'hbce68529; // ẋ171:-0.028139667585492134
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'hb8454a62; // θ171:-4.703773447545245e-05
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'hbbca80c0; // ω171:-0.006179898977279663

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'hbc2df212; // x172:-0.010616796091198921
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'hbaefe70e; // ẋ172:-0.0018303112592548132
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h3ca2b572; // θ172:0.019861910492181778
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'hbd090cfc; // ω172:-0.03345964848995209

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h3c0eba4d; // x173:0.008711409755051136
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h3cff6ef4; // ẋ173:0.031180836260318756
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h3d36b7ad; // θ173:0.04460876062512398
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'hbca34f26; // ω173:-0.019935201853513718

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'hbce1cf36; // x174:-0.027564626187086105
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'hbad2adcb; // ẋ174:-0.0016073522856459022
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h3d4adf85; // θ174:0.04952957108616829
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h3d416b5d; // ω174:0.047221530228853226

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'hbc9c5192; // x175:-0.01908186450600624
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'hbb6c1b88; // ẋ175:-0.0036027152091264725
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'hbd306064; // θ175:-0.043060675263404846
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h3c2e33aa; // ω175:0.010632434859871864

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'hbcef311e; // x176:-0.02919822558760643
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'hbd3ff7d2; // ẋ176:-0.04686719924211502
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'hbd207572; // θ176:-0.039174504578113556
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h3d1a5209; // ω176:0.037675891071558

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'hbc409685; // x177:-0.011754636652767658
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h3d1bb3eb; // ẋ177:0.03801338002085686
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'hbd471bf8; // θ177:-0.04861065745353699
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'hbba8d0df; // ω177:-0.005151852499693632

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'hbd121f03; // x178:-0.03567410632967949
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'hbbb605c1; // ẋ178:-0.005554885137826204
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'hbd49602a; // θ178:-0.049163974821567535
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h3d21e3c3; // ω178:0.03952385112643242

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h3d0d4061; // x179:0.03448522463440895
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'hbabbce7b; // ẋ179:-0.0014328503748402
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'hbca06d3b; // θ179:-0.019583335146307945
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'hbd2e034d; // ω179:-0.0424836166203022

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'hbc8b7f6b; // x180:-0.017028531059622765
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'hbd4a4536; // ẋ180:-0.04938241094350815
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h3cc6120d; // θ180:0.024178529158234596
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h3cea3323; // ω180:0.028588837012648582

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'hbc91de7a; // x181:-0.0178062804043293
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'hbd24a71c; // ẋ181:-0.0401984304189682
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'hbd0407ad; // θ181:-0.03223388269543648
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'hbcd3adc0; // ω181:-0.025839686393737793

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'hbd4b0ca1; // x182:-0.04957259073853493
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h3d3fdcca; // ẋ182:0.046841420233249664
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h3d461ecd; // θ182:0.04836921766400337
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h3ceb8454; // ω182:0.028749622404575348

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h3c6164ad; // x183:0.013756913132965565
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h3b602b33; // ẋ183:0.003420543624088168
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h3d2071f8; // θ183:0.039171189069747925
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h3d0fb926; // ω183:0.0350886806845665

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h3c139ced; // x184:0.009009581990540028
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h3d2cc6c5; // ẋ184:0.042181748896837234
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h3cef1368; // θ184:0.02918405830860138
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h3d266a4b; // ω184:0.04062871262431145

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'hbc86f102; // x185:-0.01647234335541725
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h3d191c30; // ẋ185:0.0373803973197937
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'hbc8b913e; // θ185:-0.017037030309438705
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'hbb22d458; // ω185:-0.0024845805019140244

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'hbd495f77; // x186:-0.04916330799460411
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h3c0f1b59; // ẋ186:0.008734547533094883
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'hb9465906; // θ186:-0.00018915915279649198
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'hbd171c41; // ω186:-0.036892179399728775

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h3ce50727; // x187:0.027957512065768242
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'hbc9af6bf; // ẋ187:-0.018916485831141472
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'hbd4c63bc; // θ187:-0.04989980161190033
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'hbd159e7b; // ω187:-0.0365280918776989

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h3cc90b10; // x188:0.024541407823562622
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'hbd157025; // ẋ188:-0.03648390248417854
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'hbcb3271d; // θ188:-0.02186923660337925
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'hbcd01e6c; // ω188:-0.02540513128042221

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'hbc1243d6; // x189:-0.008927306160330772
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'hbcef841d; // ẋ189:-0.02923780120909214
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h3d493d46; // θ189:0.049130700528621674
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'hbd25c0aa; // ω189:-0.04046694189310074

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'hbabec383; // x190:-0.00145541166421026
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h3cbbfac9; // ẋ190:0.022946732118725777
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'hbc8fcb07; // θ190:-0.01755286566913128
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h3cace5af; // ω190:0.02110561542212963

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'hbcf268ea; // x191:-0.029591042548418045
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'hbcc63671; // ẋ191:-0.024195881560444832
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'hbc1a4c37; // θ191:-0.009417585097253323
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'hbd0c5d8a; // ω191:-0.03426889330148697

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'hbd1fdd0b; // x192:-0.039029162377119064
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h3d238d8f; // ẋ192:0.03992992267012596
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h3c7e216c; // θ192:0.01551089808344841
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'hbc8200aa; // ω192:-0.01586945727467537

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h3d2612b3; // x193:0.04054517671465874
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'hbd21b660; // ẋ193:-0.03948056697845459
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h3c335b25; // θ193:0.010947023518383503
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'hbd0b6c66; // ω193:-0.03403892368078232

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'hbd01ae99; // x194:-0.03166064992547035
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'hbc7233cb; // ẋ194:-0.014782856218516827
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'hbd4253d4; // θ194:-0.04744322597980499
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h3cb35f3a; // ω194:0.021895993500947952

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h3d4a7690; // x195:0.049429476261138916
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h3c97c93a; // ẋ195:0.018528569489717484
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h3d124205; // θ195:0.035707492381334305
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h3d18c74f; // ω195:0.03729945048689842

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h3c474039; // x196:0.012161307968199253
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h3b7fa5b6; // ẋ196:0.0039008683525025845
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h3c2e0ef0; // θ196:0.01062367856502533
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'hbc9802b4; // ω196:-0.018555976450443268

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'hbb07bc7e; // x197:-0.002071171533316374
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h3d3b898d; // ẋ197:0.04578547552227974
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'hbd272ca5; // θ197:-0.04081406071782112
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h3cb1afd2; // ω197:0.021690282970666885

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'hbcfc23a4; // x198:-0.030778713524341583
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h3cfb4ced; // ẋ198:0.030676329508423805
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'hbcceec22; // θ198:-0.02525908127427101
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'hbd29cd3f; // ω198:-0.041455503553152084

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'hbcaf3014; // x199:-0.021385230123996735
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h3cd886fb; // ẋ199:0.026431551203131676
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'hbd3a70a7; // θ199:-0.04551758989691734
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'hbd182c39; // ω199:-0.03715154901146889

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h3c938fce; // x200:0.01801290735602379
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h3d43c8bf; // ẋ200:0.047798868268728256
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h3d4602fb; // θ200:0.048342686146497726
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'hbc50d174; // ω200:-0.012745250016450882

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h3cdc9fb8; // x201:0.026931628584861755
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'hbcce174b; // ẋ201:-0.025157591328024864
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h3d3a6f70; // θ201:0.04551643133163452
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'hbb35323c; // ω201:-0.0027648350223898888

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'hbd1fb50b; // x202:-0.038991015404462814
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h3b87c0d0; // ẋ202:0.00414285808801651
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'hbce82d7c; // θ202:-0.028342001140117645
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'hbce79dd4; // ω202:-0.028273500502109528

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'hbcf10c26; // x203:-0.02942473813891411
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h3c4e0b1e; // ẋ203:0.012575892731547356
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'hbd46d57e; // θ203:-0.04854344576597214
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h3d1dd8d9; // ω203:0.038536880165338516

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'hbbbad90b; // x204:-0.00570214306935668
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h3cbd41d8; // ẋ204:0.023102685809135437
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h3cdb7e1e; // θ204:0.02679353579878807
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'hbd1e2e32; // ω204:-0.03861827403306961

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h3c2f0556; // x205:0.010682424530386925
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'hbccf8959; // ẋ205:-0.02533404715359211
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h3c518a06; // θ205:0.012789255008101463
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h3bc3d39c; // ω205:0.005976153537631035

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h3c9a704f; // x206:0.01885238103568554
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h3d399869; // ẋ206:0.04531136527657509
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'hbd3fae96; // θ206:-0.04679735749959946
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h3c04ed76; // ω206:0.008113255724310875

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'hbb92844d; // x207:-0.004471337888389826
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h3ad1772d; // ẋ207:0.001598095172084868
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h3d14bccd; // θ207:0.03631286695599556
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'hbcc91e7a; // ω207:-0.0245506651699543

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h3d4c920c; // x208:0.049943968653678894
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h3d329c50; // ẋ208:0.04360610246658325
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'hbbfe4b47; // θ208:-0.0077604386024177074
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h3ccb89cf; // ω208:0.02484598569571972

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'hbccc7226; // x209:-0.024956773966550827
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h3d1e3158; // ẋ209:0.03862127661705017
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'hbb90b1db; // θ209:-0.004415733274072409
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'hba44dd94; // ω209:-0.0007509824354201555

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'hbd010261; // x210:-0.03149640932679176
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h3ce9d599; // ẋ210:0.028544234111905098
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h3c95219f; // θ210:0.01820450834929943
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'hbbe127bf; // ω210:-0.006871193181723356

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h3c9b1bb9; // x211:0.018934117630124092
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'hba330b0a; // ẋ211:-0.0006829953053966165
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h3d0931da; // θ211:0.03349480777978897
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'hbc8a424e; // ω211:-0.016877319663763046

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h3c15232f; // x212:0.009102626703679562
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h3c2415c7; // ẋ212:0.010014957748353481
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h3d3ba149; // θ212:0.045808110386133194
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'hbc2be2a1; // ω212:-0.010491044260561466

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'hbc6777ea; // x213:-0.014127710834145546
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'hbcbafb06; // ẋ213:-0.02282477542757988
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'hbcb9f407; // θ213:-0.022699369117617607
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h3cf977bb; // ω213:0.030452599748969078

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'hbb007322; // x214:-0.001959987450391054
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'hba49c783; // ẋ214:-0.0007697271066717803
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'hbcc0c493; // θ214:-0.02353123389184475
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'hbc7a28f5; // ω214:-0.015268553979694843

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h3c9198e1; // x215:0.017773093655705452
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'hbd42074d; // ẋ215:-0.047370243817567825
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'hbab8976a; // θ215:-0.0014083210844546556
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'hbca07ace; // ω215:-0.019589807838201523

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h3d0ec389; // x216:0.03485444560647011
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h3ca80ab0; // ẋ216:0.020512908697128296
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'hbd0c6977; // θ216:-0.03428026661276817
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h3c98f414; // ω216:0.018671073019504547

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h3cdbd6ce; // x217:0.02683582529425621
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'hbbc1a5d7; // ẋ217:-0.00590966222807765
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'hbd041dd7; // θ217:-0.03225501999258995
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h3cee4412; // ω217:0.0290851928293705

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'hbd282d51; // x218:-0.04105884209275246
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h3bdd1652; // ẋ218:0.006747045554220676
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'hbd3148a2; // θ218:-0.0432821586728096
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h3d06cf42; // ω218:0.03291250020265579

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'hbc49fb2d; // x219:-0.01232795137912035
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'hbc8df6a1; // ẋ219:-0.017329515889286995
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h3bcb5e4d; // θ219:0.006206309888511896
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h3cbf4850; // ω219:0.023349910974502563

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h3d42c449; // x220:0.04755047336220741
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'hbd2e500a; // ẋ220:-0.042556799948215485
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'hbc6bb752; // θ220:-0.014386968687176704
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h3cb07ba7; // ω220:0.021543337032198906

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'hbd2e9955; // x221:-0.042626697570085526
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'hbbdb7eeb; // ẋ221:-0.006698479410260916
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h3b187902; // θ221:0.0023265485651791096
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h3d3e3dc2; // ω221:0.04644561558961868

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'hbd43e5e5; // x222:-0.04782666638493538
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h3c28fe15; // ẋ222:0.010314484126865864
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h3cf183c6; // θ222:0.029481779783964157
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h3b626045; // ω222:0.0034542244393378496

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h3c2e51a3; // x223:0.010639580897986889
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'hbd2a2905; // ẋ223:-0.04154302552342415
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h3b957d86; // θ223:0.004562082700431347
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h3d2b5788; // ω223:0.041831523180007935

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h3ca51221; // x224:0.02015024609863758
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h3c2253eb; // ẋ224:0.009907702915370464
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h3c9f4eac; // θ224:0.01944669336080551
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'hbc05c3fe; // ω224:-0.008164403960108757

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'hbbc600ad; // x225:-0.006042561028152704
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'hbca30b1e; // ẋ225:-0.01990276202559471
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h3ce1d800; // θ225:0.027568817138671875
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'hbd12d61d; // ω225:-0.03584872558712959

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'hbd0474c7; // x226:-0.03233793005347252
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'hbc828d7f; // ẋ226:-0.015936611220240593
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h3a8f3ed5; // θ226:0.0010928759584203362
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h3cbca9f4; // ω226:0.02303025871515274

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h3cc24593; // x227:0.023714816197752953
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'hbb0ddeb6; // ẋ227:-0.0021647638641297817
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h3cce9a29; // θ227:0.0252199936658144
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'hbbd625e2; // ω227:-0.0065352777019143105

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h3c337dfa; // x228:0.01095532812178135
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h3d43febf; // ẋ228:0.047850366681814194
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'hbc9a6b41; // θ228:-0.018849970772862434
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'hbcd2400b; // ω228:-0.02566530369222164

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h3c87d39f; // x229:0.016580400988459587
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'hbc500bd1; // ẋ229:-0.012698129750788212
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h3bb8bc75; // θ229:0.005637700203806162
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'hbca8b62e; // ω229:-0.020594682544469833

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h3d0635e0; // x230:0.03276622295379639
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'hbd1da2cc; // ẋ230:-0.0384853333234787
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'hbc0e033a; // θ230:-0.008667761459946632
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h3c6e0918; // ω230:0.014528535306453705

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'hbd3d6dfa; // x231:-0.0462474599480629
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'hbd31e62c; // ẋ231:-0.04343239963054657
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h3cd29142; // θ231:0.025704029947519302
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'hbd01379a; // ω231:-0.03154716640710831

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'hbd10edfc; // x232:-0.035383209586143494
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h3be5ad1a; // ẋ232:0.007009160704910755
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h3cfdf728; // θ232:0.03100164234638214
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'hbd28a4b2; // ω232:-0.04117269068956375

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'hbb82967c; // x233:-0.003985224291682243
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'hbd217805; // ẋ233:-0.03942110016942024
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h3cd15557; // θ233:0.02555338852107525
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'hb7b48831; // ω233:-2.152109118469525e-05

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'hbcd2ace9; // x234:-0.02571721561253071
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h3d36c43f; // ẋ234:0.04462074860930443
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'hbcf78379; // θ234:-0.030214058235287666
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'hbb3b515a; // ω234:-0.0028582424856722355

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'hbcb4d2c4; // x235:-0.022073157131671906
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'hbcc94824; // ẋ235:-0.024570532143115997
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'hbba8b27a; // θ235:-0.005148229189217091
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h3c8424ec; // ω235:0.01613088697195053

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'hbd15f767; // x236:-0.036612894386053085
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h3d1a5bc1; // ẋ236:0.03768515959382057
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h3d064739; // θ236:0.032782766968011856
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h3c806431; // ω236:0.015672774985432625

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h3aacbdb0; // x237:0.001317908987402916
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'hbc99d576; // ẋ237:-0.018778543919324875
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'hbd2f3715; // θ237:-0.04277713969349861
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h39de6a72; // ω237:0.000424224475864321

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h3a57ee7b; // x238:0.0008237135480158031
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h3cb4192b; // ẋ238:0.021984657272696495
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h3c9efb1c; // θ238:0.019406847655773163
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h3b4f33d3; // ω238:0.003161658300086856

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'hbd48dc20; // x239:-0.049038052558898926
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h3c1975a0; // ẋ239:0.009366422891616821
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'hbcb053ef; // θ239:-0.021524397656321526
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h3b1295f4; // ω239:0.0022367211058735847

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'hbd000191; // x240:-0.03125149384140968
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'h3c01292e; // ẋ240:0.007883353158831596
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'h3cd4ef52; // θ240:0.025993023067712784
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'hbca57b71; // ω240:-0.020200463011860847

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'h3ba243fa; // x241:0.004951951093971729
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'h3d1cdcc7; // ẋ241:0.03829648718237877
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'hbb790aaa; // θ241:-0.003800074104219675
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd967; ram_i_data1 = 32'h3d000f57; // ω241:0.03126462921500206

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd968; ram_i_data1 = 32'h3c247108; // x242:0.010036714375019073
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd969; ram_i_data1 = 32'hbb168f3e; // ẋ242:-0.0022973562590777874
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd970; ram_i_data1 = 32'hbb8555fd; // θ242:-0.004069088492542505
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd971; ram_i_data1 = 32'hbd3a533b; // ω242:-0.04548953101038933

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd972; ram_i_data1 = 32'hbccf748e; // x243:-0.025324132293462753
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd973; ram_i_data1 = 32'h3d03ab13; // ẋ243:0.03214557096362114
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd974; ram_i_data1 = 32'hbd426901; // θ243:-0.047463420778512955
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd975; ram_i_data1 = 32'hbd3714d5; // ω243:-0.0446976013481617

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd976; ram_i_data1 = 32'h3d43d921; // x244:0.047814492136240005
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd977; ram_i_data1 = 32'h3d167ade; // ẋ244:0.03673826903104782
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd978; ram_i_data1 = 32'hbc435ef1; // θ244:-0.01192449126392603
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd979; ram_i_data1 = 32'h3d1508a4; // ω244:0.0363851934671402

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd980; ram_i_data1 = 32'hbd27fce3; // x245:-0.041012655943632126
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd981; ram_i_data1 = 32'hbb8a4d6e; // ẋ245:-0.004220656119287014
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd982; ram_i_data1 = 32'h3ce391f9; // θ245:0.02777956612408161
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd983; ram_i_data1 = 32'h3b6caf8a; // ω245:0.0036115371622145176

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd984; ram_i_data1 = 32'hbd3003f4; // x246:-0.04297251999378204
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd985; ram_i_data1 = 32'hbc2138f1; // ẋ246:-0.00984023604542017
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd986; ram_i_data1 = 32'h3c3e6f06; // θ246:0.011623149737715721
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd987; ram_i_data1 = 32'hbd303859; // ω246:-0.04302248731255531

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd988; ram_i_data1 = 32'hbd214bb4; // x247:-0.03937883675098419
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd989; ram_i_data1 = 32'h3d113d43; // ẋ247:0.03545881435275078
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd990; ram_i_data1 = 32'hbcaf94bd; // θ247:-0.021433228626847267
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd991; ram_i_data1 = 32'h3d191399; // ω247:0.03737220540642738

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd992; ram_i_data1 = 32'hbc87e248; // x248:-0.01658739149570465
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd993; ram_i_data1 = 32'h3d3df85d; // ẋ248:0.04637943580746651
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd994; ram_i_data1 = 32'h3c87ebea; // θ248:0.016591984778642654
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd995; ram_i_data1 = 32'hbd24bffe; // ω248:-0.0402221605181694

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd996; ram_i_data1 = 32'hbd4160b6; // x249:-0.04721137136220932
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd997; ram_i_data1 = 32'h3c8ee7b7; // ẋ249:0.01744447462260723
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd998; ram_i_data1 = 32'h3cb36fd7; // θ249:0.02190391533076763
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd999; ram_i_data1 = 32'hbc524a58; // ω249:-0.012835107743740082

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1000; ram_i_data1 = 32'hbcf04ab3; // x250:-0.029332494363188744
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1001; ram_i_data1 = 32'h3b88ee1c; // ẋ250:0.0041787754744291306
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1002; ram_i_data1 = 32'hbc1a782e; // θ250:-0.00942806713283062
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1003; ram_i_data1 = 32'h3ba78e8b; // ω250:0.005113427992910147

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1004; ram_i_data1 = 32'h3ba16a42; // x251:0.004925996996462345
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1005; ram_i_data1 = 32'h3b2b61eb; // ẋ251:0.0026150892954319715
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1006; ram_i_data1 = 32'hbc5bdb31; // θ251:-0.013418958522379398
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1007; ram_i_data1 = 32'h3d3d382e; // ω251:0.04619615525007248

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1008; ram_i_data1 = 32'h3d1dc0ba; // x252:0.038513876497745514
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1009; ram_i_data1 = 32'hbce242e6; // ẋ252:-0.02761979028582573
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1010; ram_i_data1 = 32'h3c9012f2; // θ252:0.01758715882897377
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1011; ram_i_data1 = 32'hbd0b8976; // ω252:-0.034066639840602875

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1012; ram_i_data1 = 32'h3d03d109; // x253:0.03218177333474159
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1013; ram_i_data1 = 32'h3cdb563b; // ẋ253:0.026774516329169273
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1014; ram_i_data1 = 32'h3bcfc9f4; // θ253:0.00634121336042881
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1015; ram_i_data1 = 32'hbd28c166; // ω253:-0.04120006412267685

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1016; ram_i_data1 = 32'hbd0af9e1; // x254:-0.03392970934510231
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1017; ram_i_data1 = 32'h3d36eff7; // ẋ254:0.044662442058324814
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1018; ram_i_data1 = 32'h3cceed3b; // θ254:0.025259604677557945
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1019; ram_i_data1 = 32'h3d09b72f; // ω254:0.03362196311354637

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1020; ram_i_data1 = 32'hbd235b84; // x255:-0.039882197976112366
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1021; ram_i_data1 = 32'hba0d6bcd; // ẋ255:-0.000539478671271354
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1022; ram_i_data1 = 32'h3c430f9e; // θ255:0.011905578896403313
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1023; ram_i_data1 = 32'h3d1ee478; // ω255:0.03879210352897644

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1024; ram_i_data1 = 32'hbb421793; // x256:-0.002961610211059451
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1025; ram_i_data1 = 32'h3ce5b87e; // ẋ256:0.028042074292898178
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1026; ram_i_data1 = 32'hba3ff23a; // θ256:-0.0007322166347876191
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1027; ram_i_data1 = 32'h3d2beaa7; // ω256:0.041971828788518906

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1028; ram_i_data1 = 32'hbbac7983; // x257:-0.005263508763164282
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1029; ram_i_data1 = 32'hbccba89d; // ẋ257:-0.024860674515366554
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1030; ram_i_data1 = 32'h3c77b909; // θ257:0.01511979941278696
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1031; ram_i_data1 = 32'hbc66f3f1; // ω257:-0.014096246100962162

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1032; ram_i_data1 = 32'h3d0015b1; // x258:0.03127068653702736
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1033; ram_i_data1 = 32'h3ce631af; // ẋ258:0.02809986285865307
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1034; ram_i_data1 = 32'hbc6cd969; // θ258:-0.014456131495535374
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1035; ram_i_data1 = 32'hbd01316e; // ω258:-0.03154128044843674

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1036; ram_i_data1 = 32'h3b2a1018; // x259:0.002594953402876854
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1037; ram_i_data1 = 32'h3d199f0c; // ẋ259:0.037505194544792175
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1038; ram_i_data1 = 32'h3caf3f1d; // θ259:0.021392399445176125
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1039; ram_i_data1 = 32'h3d1de8fb; // ω259:0.038552265614271164

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1040; ram_i_data1 = 32'hbd24cbea; // x260:-0.04023353010416031
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1041; ram_i_data1 = 32'h3b1281d2; // ẋ260:0.0022355210967361927
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1042; ram_i_data1 = 32'hbcc7f908; // θ260:-0.024410739541053772
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1043; ram_i_data1 = 32'hbbf199aa; // ω260:-0.007373054511845112

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1044; ram_i_data1 = 32'h3d0a5d81; // x261:0.03378057852387428
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1045; ram_i_data1 = 32'hbd3b2d2c; // ẋ261:-0.045697376132011414
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1046; ram_i_data1 = 32'hbd43944e; // θ261:-0.047748856246471405
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1047; ram_i_data1 = 32'hbc77da7a; // ω261:-0.015127772465348244

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1048; ram_i_data1 = 32'h3d2977c8; // x262:0.041373997926712036
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1049; ram_i_data1 = 32'hba6d5f72; // ẋ262:-0.0009055054979398847
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1050; ram_i_data1 = 32'hbc3c9245; // θ262:-0.011509482748806477
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1051; ram_i_data1 = 32'hbd42f937; // ω262:-0.04760095104575157

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1052; ram_i_data1 = 32'hbbae5463; // x263:-0.005320118274539709
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1053; ram_i_data1 = 32'hbcda20b9; // ẋ263:-0.026626931503415108
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1054; ram_i_data1 = 32'h3cf130b0; // θ263:0.029442161321640015
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1055; ram_i_data1 = 32'h3bc04b44; // ω263:0.0058683473616838455

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1056; ram_i_data1 = 32'hbce4f5af; // x264:-0.02794918231666088
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1057; ram_i_data1 = 32'h3d47099a; // ẋ264:0.04859314113855362
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1058; ram_i_data1 = 32'hbd22d26c; // θ264:-0.039751455187797546
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1059; ram_i_data1 = 32'hbbda27e1; // ω264:-0.006657585967332125

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1060; ram_i_data1 = 32'h3d16a4ef; // x265:0.03677838668227196
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1061; ram_i_data1 = 32'hbca1c67a; // ẋ265:-0.019747961312532425
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1062; ram_i_data1 = 32'hbd482ce0; // θ265:-0.04887092113494873
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1063; ram_i_data1 = 32'hba5a2652; // ω265:-0.0008321750210598111

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1064; ram_i_data1 = 32'hbc394250; // x266:-0.011307314038276672
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1065; ram_i_data1 = 32'hbc0ad964; // ẋ266:-0.0084746815264225
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1066; ram_i_data1 = 32'h3d1c4a60; // θ266:0.038156867027282715
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1067; ram_i_data1 = 32'hbd1f408c; // ω266:-0.038879916071891785

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1068; ram_i_data1 = 32'hbb65a6f5; // x267:-0.00350421410985291
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1069; ram_i_data1 = 32'hbd303889; // ẋ267:-0.04302266612648964
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1070; ram_i_data1 = 32'hbd456a5a; // θ267:-0.048197127878665924
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1071; ram_i_data1 = 32'h3c87ec52; // ω267:0.016592178493738174

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1072; ram_i_data1 = 32'h3d064e2c; // x268:0.03278939425945282
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1073; ram_i_data1 = 32'h3d3d58e9; // ẋ268:0.04622736945748329
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1074; ram_i_data1 = 32'h3c0acbe1; // θ268:0.008471460081636906
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1075; ram_i_data1 = 32'h3cf8aff5; // ω268:0.03035734035074711

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1076; ram_i_data1 = 32'h3d380f40; // x269:0.044936418533325195
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1077; ram_i_data1 = 32'hbd3b8b43; // ẋ269:-0.045787107199430466
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1078; ram_i_data1 = 32'h3c912bae; // θ269:0.0177210234105587
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1079; ram_i_data1 = 32'hbcced88a; // ω269:-0.02524973824620247

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1080; ram_i_data1 = 32'h3d1d44d8; // x270:0.03839573264122009
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1081; ram_i_data1 = 32'hbc2cfcd2; // ẋ270:-0.010558323934674263
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1082; ram_i_data1 = 32'hbc25d457; // θ270:-0.010121426545083523
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1083; ram_i_data1 = 32'hbd0cb894; // ω270:-0.03435571491718292

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1084; ram_i_data1 = 32'h3d073717; // x271:0.03301152214407921
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1085; ram_i_data1 = 32'h3ccd234a; // ẋ271:0.025041241198778152
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1086; ram_i_data1 = 32'hbd3db2b6; // θ271:-0.04631301015615463
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1087; ram_i_data1 = 32'hbcd1e65c; // ω271:-0.025622539222240448

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1088; ram_i_data1 = 32'h3cbb7fdc; // x272:0.022888116538524628
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1089; ram_i_data1 = 32'hbd36fa88; // ẋ272:-0.04467251896858215
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1090; ram_i_data1 = 32'hbb143cda; // θ272:-0.00226192781701684
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1091; ram_i_data1 = 32'hbc81e70b; // ω272:-0.015857240185141563

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1092; ram_i_data1 = 32'hbd2f139a; // x273:-0.04274330288171768
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1093; ram_i_data1 = 32'hbab8ea7c; // ẋ273:-0.0014107967726886272
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1094; ram_i_data1 = 32'hbc169948; // θ273:-0.009191818535327911
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1095; ram_i_data1 = 32'hbc0168bd; // ω273:-0.007898506708443165

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1096; ram_i_data1 = 32'hbcc08783; // x274:-0.02350211702287197
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1097; ram_i_data1 = 32'h3c22ab77; // ẋ274:0.009928575716912746
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1098; ram_i_data1 = 32'hbc3d5db1; // θ274:-0.011557982303202152
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1099; ram_i_data1 = 32'hbd3043db; // ω274:-0.04303346201777458

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1100; ram_i_data1 = 32'h3b4572db; // x275:0.0030128273647278547
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1101; ram_i_data1 = 32'h3c8c13d9; // ẋ275:0.017099307850003242
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1102; ram_i_data1 = 32'hbd4147ff; // θ275:-0.04718780145049095
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1103; ram_i_data1 = 32'h3c4f5d0c; // ω275:0.01265646144747734

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1104; ram_i_data1 = 32'h3a1260e9; // x276:0.0005583898746408522
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1105; ram_i_data1 = 32'h3d036a51; // ẋ276:0.03208381310105324
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1106; ram_i_data1 = 32'hbc7bf93a; // θ276:-0.015379244461655617
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1107; ram_i_data1 = 32'hbcf02848; // ω276:-0.02931608259677887

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1108; ram_i_data1 = 32'h3aec5dba; // x277:0.0018033303786069155
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1109; ram_i_data1 = 32'hbc01b00f; // ẋ277:-0.007915510796010494
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1110; ram_i_data1 = 32'hbbe4adf9; // θ277:-0.006978746969252825
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1111; ram_i_data1 = 32'hbd3cbf99; // ω277:-0.04608115926384926

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1112; ram_i_data1 = 32'h3c0309cd; // x278:0.00799794215708971
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1113; ram_i_data1 = 32'h3cae1873; // ẋ278:0.021251892670989037
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1114; ram_i_data1 = 32'hbd1b9ee3; // θ278:-0.03799332305788994
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1115; ram_i_data1 = 32'hbd16a764; // ω278:-0.03678072988986969

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1116; ram_i_data1 = 32'h3ca04b2c; // x279:0.0195670947432518
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1117; ram_i_data1 = 32'hbce9dc4f; // ẋ279:-0.028547434136271477
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1118; ram_i_data1 = 32'h3c015fd4; // θ279:0.007896382361650467
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1119; ram_i_data1 = 32'hbca25488; // ω279:-0.019815698266029358

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1120; ram_i_data1 = 32'h3d12eff2; // x280:0.03587336093187332
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1121; ram_i_data1 = 32'h3d41defc; // ẋ280:0.0473317950963974
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1122; ram_i_data1 = 32'hbca056a1; // θ280:-0.019572557881474495
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1123; ram_i_data1 = 32'h3cb32eab; // ω280:0.021872838959097862

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1124; ram_i_data1 = 32'hbcb41051; // x281:-0.021980436518788338
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1125; ram_i_data1 = 32'hbd168711; // ẋ281:-0.03674990311264992
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1126; ram_i_data1 = 32'h3cf0d953; // θ281:0.029400503262877464
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1127; ram_i_data1 = 32'hbd2cc1fe; // ω281:-0.042177192866802216

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1128; ram_i_data1 = 32'h3c82c561; // x282:0.01596325822174549
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1129; ram_i_data1 = 32'hbc8767b3; // ẋ282:-0.016528939828276634
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1130; ram_i_data1 = 32'hbd40c94b; // θ282:-0.04706696793437004
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1131; ram_i_data1 = 32'h3cf86ae1; // ω282:0.030324401333928108

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1132; ram_i_data1 = 32'h3d02bd14; // x283:0.03191860020160675
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1133; ram_i_data1 = 32'hbd4587b4; // ẋ283:-0.04822511970996857
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1134; ram_i_data1 = 32'hbc48cd89; // θ283:-0.012256034649908543
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1135; ram_i_data1 = 32'hbaf7ef41; // ω283:-0.001891590771265328

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1136; ram_i_data1 = 32'hbd171418; // x284:-0.03688439726829529
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1137; ram_i_data1 = 32'hbb6dcd73; // ẋ284:-0.0036285787355154753
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1138; ram_i_data1 = 32'h3d2d9f56; // θ284:0.04238828271627426
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1139; ram_i_data1 = 32'h3d32ab8b; // ω284:0.043620627373456955

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1140; ram_i_data1 = 32'hbb983177; // x285:-0.004644568543881178
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1141; ram_i_data1 = 32'h3ce6415a; // ẋ285:0.028107333928346634
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1142; ram_i_data1 = 32'hbcb25685; // θ285:-0.021769771352410316
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1143; ram_i_data1 = 32'h3cf00b98; // ω285:0.029302403330802917

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1144; ram_i_data1 = 32'hbca5e773; // x286:-0.020251965150237083
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1145; ram_i_data1 = 32'hbd421cce; // ẋ286:-0.04739075154066086
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1146; ram_i_data1 = 32'hba9cd083; // θ286:-0.0011963996803388
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1147; ram_i_data1 = 32'hbd3ec764; // ω286:-0.04657687246799469

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1148; ram_i_data1 = 32'h3c111031; // x287:0.008853957988321781
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1149; ram_i_data1 = 32'hbb80a7e0; // ẋ287:-0.003926262259483337
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1150; ram_i_data1 = 32'hbc92dc4b; // θ287:-0.01792730949819088
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1151; ram_i_data1 = 32'hbcd37a60; // ω287:-0.025815188884735107

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1152; ram_i_data1 = 32'h3d0fac68; // x288:0.035076528787612915
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1153; ram_i_data1 = 32'h3cdf3e69; // ẋ288:0.027251439169049263
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1154; ram_i_data1 = 32'hbc26b77b; // θ288:-0.010175581090152264
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1155; ram_i_data1 = 32'h3d237682; // ω288:0.03990793973207474

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1156; ram_i_data1 = 32'h3ba837bb; // x289:0.0051335967145860195
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1157; ram_i_data1 = 32'h3d191486; // ẋ289:0.03737308830022812
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1158; ram_i_data1 = 32'h3ce47022; // θ289:0.027885500341653824
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1159; ram_i_data1 = 32'h3d0098a1; // ω289:0.0313955582678318

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1160; ram_i_data1 = 32'hbcd326e0; // x290:-0.025775372982025146
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1161; ram_i_data1 = 32'hbd4c7330; // ẋ290:-0.049914538860321045
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1162; ram_i_data1 = 32'h3d06bcbe; // θ290:0.03289484232664108
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1163; ram_i_data1 = 32'hbb76b62e; // ω290:-0.003764520864933729

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1164; ram_i_data1 = 32'h3cd8b383; // x291:0.02645278535783291
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1165; ram_i_data1 = 32'hbca22616; // ẋ291:-0.019793551415205002
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1166; ram_i_data1 = 32'h3d42f834; // θ291:0.04759998619556427
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1167; ram_i_data1 = 32'h3d14cffb; // ω291:0.03633115813136101

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1168; ram_i_data1 = 32'h3c2c2c3f; // x292:0.01050859596580267
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1169; ram_i_data1 = 32'h3d090dc1; // ẋ292:0.033460382372140884
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1170; ram_i_data1 = 32'hbcf57a9b; // θ292:-0.029965689405798912
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1171; ram_i_data1 = 32'h3a7b6902; // ω292:0.0009590537520125508

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1172; ram_i_data1 = 32'h3cda4d63; // x293:0.026648228988051414
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1173; ram_i_data1 = 32'hbcff1bab; // ẋ293:-0.031141122803092003
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1174; ram_i_data1 = 32'hbcd694ec; // θ293:-0.02619405835866928
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1175; ram_i_data1 = 32'hbd1dde98; // ω293:-0.038542360067367554

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1176; ram_i_data1 = 32'hbc28d8c4; // x294:-0.010305587202310562
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1177; ram_i_data1 = 32'h3c793560; // ẋ294:0.015210479497909546
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1178; ram_i_data1 = 32'h3bbe1761; // θ294:0.005801126826554537
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1179; ram_i_data1 = 32'hbd09c64d; // ω294:-0.03363637998700142

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1180; ram_i_data1 = 32'hbca9c84d; // x295:-0.020725393667817116
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1181; ram_i_data1 = 32'hbccba33a; // ẋ295:-0.024858105927705765
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1182; ram_i_data1 = 32'h3d2e9137; // θ295:0.04261895641684532
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1183; ram_i_data1 = 32'hbc9c77db; // ω295:-0.019100120291113853

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1184; ram_i_data1 = 32'h3d216819; // x296:0.03940591588616371
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1185; ram_i_data1 = 32'hbba1ce81; // ẋ296:-0.004937947262078524
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1186; ram_i_data1 = 32'hbd0f1a95; // θ296:-0.03493745997548103
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1187; ram_i_data1 = 32'hbb333a52; // ω296:-0.0027347994036972523

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1188; ram_i_data1 = 32'hbc436307; // x297:-0.011925465427339077
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1189; ram_i_data1 = 32'hbb592f42; // ẋ297:-0.0033139740116894245
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1190; ram_i_data1 = 32'hbad9a60e; // θ297:-0.001660527428612113
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1191; ram_i_data1 = 32'h3d07f68d; // ω297:0.03319411352276802

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1192; ram_i_data1 = 32'hbbf59711; // x298:-0.007494815159589052
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1193; ram_i_data1 = 32'h3ca5ce35; // ẋ298:0.020239928737282753
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1194; ram_i_data1 = 32'h3d3670c6; // θ298:0.044541142880916595
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1195; ram_i_data1 = 32'h3cd83644; // ω298:0.026393063366413116

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1196; ram_i_data1 = 32'hbcc2fd53; // x299:-0.023802435025572777
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1197; ram_i_data1 = 32'h3c14b3ab; // ẋ299:0.009076039306819439
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1198; ram_i_data1 = 32'h3cf84262; // θ299:0.03030509129166603
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1199; ram_i_data1 = 32'hbc5944a6; // ω299:-0.013260995969176292

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1200; ram_i_data1 = 32'hbba620a1; // x300:-0.0050698076374828815
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1201; ram_i_data1 = 32'hbd0023c6; // ẋ300:-0.031284116208553314
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1202; ram_i_data1 = 32'hbd2479a3; // θ300:-0.040155064314603806
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1203; ram_i_data1 = 32'h3ce5200d; // ω300:0.02796938456594944

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1204; ram_i_data1 = 32'h3d0e2739; // x301:0.034705374389886856
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1205; ram_i_data1 = 32'hbd26e7bc; // ẋ301:-0.040748342871665955
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1206; ram_i_data1 = 32'h3cd50618; // θ301:0.0260038822889328
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1207; ram_i_data1 = 32'h3d0faf75; // ω301:0.035079438239336014

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1208; ram_i_data1 = 32'hbd29825a; // x302:-0.041384078562259674
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1209; ram_i_data1 = 32'hbd3cf25c; // ẋ302:-0.04612956941127777
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1210; ram_i_data1 = 32'hbc083455; // θ302:-0.008313258178532124
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1211; ram_i_data1 = 32'h3d03165c; // ω302:0.032003745436668396

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1212; ram_i_data1 = 32'hbb9252c5; // x303:-0.004465433303266764
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1213; ram_i_data1 = 32'hbcfda3e4; // ẋ303:-0.030961938202381134
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1214; ram_i_data1 = 32'hbc9bd982; // θ303:-0.019024614244699478
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1215; ram_i_data1 = 32'hbc7f00f9; // ω303:-0.01556419674307108

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1216; ram_i_data1 = 32'hbd2ceccd; // x304:-0.04221801832318306
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1217; ram_i_data1 = 32'h3d4014e2; // ẋ304:0.04689491540193558
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1218; ram_i_data1 = 32'h3d2992a9; // θ304:0.04139963164925575
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1219; ram_i_data1 = 32'h3bd7843d; // ω304:0.006577043328434229

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1220; ram_i_data1 = 32'hbd18a267; // x305:-0.037264253944158554
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1221; ram_i_data1 = 32'h3d19b297; // ẋ305:0.03752383217215538
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1222; ram_i_data1 = 32'hbc9f2647; // θ305:-0.019427431747317314
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1223; ram_i_data1 = 32'h3d091301; // ω305:0.03346538916230202

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1224; ram_i_data1 = 32'hbd4b50e1; // x306:-0.049637679010629654
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1225; ram_i_data1 = 32'hbb94dce0; // ẋ306:-0.004542931914329529
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1226; ram_i_data1 = 32'hbce22537; // θ306:-0.027605636045336723
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1227; ram_i_data1 = 32'h3c3c9d52; // ω306:0.011512117460370064

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1228; ram_i_data1 = 32'h3a9a444b; // x307:0.0011769620468840003
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1229; ram_i_data1 = 32'hbd467df3; // ẋ307:-0.04845995828509331
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1230; ram_i_data1 = 32'hbc8ae6b0; // θ307:-0.016955703496932983
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1231; ram_i_data1 = 32'hbbd773c4; // ω307:-0.006575079634785652

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1232; ram_i_data1 = 32'hbcade0bc; // x308:-0.021225325763225555
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1233; ram_i_data1 = 32'h3bcbd42a; // ẋ308:0.0062203602865338326
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1234; ram_i_data1 = 32'hbce5798a; // θ308:-0.028012055903673172
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1235; ram_i_data1 = 32'hbd385512; // ω308:-0.045003004372119904

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1236; ram_i_data1 = 32'h3d3830bd; // x309:0.04496835544705391
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1237; ram_i_data1 = 32'h3d4a3fa5; // ẋ309:0.04937710240483284
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1238; ram_i_data1 = 32'h3d228126; // θ309:0.03967394679784775
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1239; ram_i_data1 = 32'h3c61a5ac; // ω309:0.013772409409284592

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1240; ram_i_data1 = 32'hbc3e4896; // x310:-0.011613985523581505
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1241; ram_i_data1 = 32'h3b346119; // ẋ310:0.0027523695025593042
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1242; ram_i_data1 = 32'h3c73eb66; // θ310:0.014887666329741478
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1243; ram_i_data1 = 32'hbcca359a; // ω310:-0.024683762341737747

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1244; ram_i_data1 = 32'h3cd76e2f; // x311:0.026297656819224358
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1245; ram_i_data1 = 32'h3d04e12d; // ẋ311:0.03244130685925484
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1246; ram_i_data1 = 32'hbd40fe6c; // θ311:-0.04711763560771942
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1247; ram_i_data1 = 32'h3d28208c; // ω311:0.041046664118766785

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1248; ram_i_data1 = 32'hbd0dd4a8; // x312:-0.03462663292884827
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1249; ram_i_data1 = 32'hbc848748; // ẋ312:-0.016177788376808167
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1250; ram_i_data1 = 32'hbd0b8792; // θ312:-0.03406483680009842
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1251; ram_i_data1 = 32'hbd0236a3; // ω312:-0.03179038688540459

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1252; ram_i_data1 = 32'hbc396dc9; // x313:-0.011317678727209568
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1253; ram_i_data1 = 32'h3d1f9125; // ẋ313:0.03895677998661995
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1254; ram_i_data1 = 32'hbd430fbe; // θ313:-0.0476224347949028
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1255; ram_i_data1 = 32'h3bd9da1a; // ω313:0.00664831418544054

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1256; ram_i_data1 = 32'h3c96a95b; // x314:0.018391301855444908
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1257; ram_i_data1 = 32'h3c4f008b; // ẋ314:0.012634406797587872
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1258; ram_i_data1 = 32'h3c2802ab; // θ314:0.010254542343318462
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1259; ram_i_data1 = 32'hbb901277; // ω314:-0.004396732430905104

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1260; ram_i_data1 = 32'h3d3cedfb; // x315:0.046125393360853195
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1261; ram_i_data1 = 32'hbcd5a12f; // ẋ315:-0.026077834889292717
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1262; ram_i_data1 = 32'hbcc1be29; // θ315:-0.023650245741009712
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1263; ram_i_data1 = 32'h3d2b3c0e; // ω315:0.04180531948804855

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1264; ram_i_data1 = 32'hbd3f9057; // x316:-0.046768512576818466
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1265; ram_i_data1 = 32'hbbfe9a72; // ẋ316:-0.007769876159727573
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1266; ram_i_data1 = 32'h3b7dc6a2; // θ316:0.0038723130710422993
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1267; ram_i_data1 = 32'hbcebc178; // ω316:-0.02877877652645111

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1268; ram_i_data1 = 32'h3d33387e; // x317:0.043755047023296356
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1269; ram_i_data1 = 32'hbc6495f6; // ẋ317:-0.013951769098639488
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1270; ram_i_data1 = 32'hbd32daee; // θ317:-0.043665818870067596
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1271; ram_i_data1 = 32'h3cec0185; // ω317:0.02880931831896305

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1272; ram_i_data1 = 32'h3c816dc6; // x318:0.01579941436648369
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1273; ram_i_data1 = 32'h3d1a9137; // ẋ318:0.03773614391684532
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1274; ram_i_data1 = 32'hbd395abc; // θ318:-0.04525254666805267
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1275; ram_i_data1 = 32'hbc3cc448; // ω318:-0.011521406471729279

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1276; ram_i_data1 = 32'hbd1d559a; // x319:-0.038411714136600494
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1277; ram_i_data1 = 32'hbc957216; // ẋ319:-0.01824287697672844
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1278; ram_i_data1 = 32'hbbd46e28; // θ319:-0.006482858210802078
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1279; ram_i_data1 = 32'hbb6e550c; // ω319:-0.003636660985648632

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 (9.0299535e26)
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.8479025e-13)
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b10101101001001110101100100001011; // action 223 ~ 192 (-9.5126225e-12)
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b11010010101011111101010111011000; // action 255 ~ 224 (-3.776035e11)
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b00100111011011000111011001110100; // action 287 ~ 256 ( 3.2815793e-15)
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b00100001101110001011000101111001; // action 319 ~ 288 ( 1.2515302e-18)

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 2nd round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b10011111100000011011111000000001; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b11100001000110000000000100110000; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b00011010110010110001100000011100; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b10011110010100000000101101001000; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b00111101101011011100010101010101; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b10011100111000001001000111110101; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b00010111011110100110000001110011; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b11000001101001001101100111110101; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b10110100110011010101000011010011; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b00010111101111101000000111101101; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 3rd round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b10011110001000100000011010100001; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b10110000010011001100100011011001; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b00011011111000110110010101110101; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b00110111011110000001111011010111; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b01001000011010001001011011000100; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b10111111110111000101110011101101; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b01010101110000100111110011111110; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b11110111101100000110000101000001; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b01010110110000111101111000001011; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b00011010110001000001111100111011; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 4th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b01010110011100001010111000101011; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b10101101101100101101101100110001; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b10111010000011001000101010100010; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b00100011011100110111101001010011; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b00101110011011001010011011011001; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b00011111101110011010011011100011; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b10111000001100011111111000000110; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b01100010000100000010000001010010; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b00101111010101100000100100100010; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b00110101011100111010101010000111; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 5th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b00011011000111001010100111111111; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b11101101001101000010001101110001; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b10100100100010010000110011101110; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b00011100011111011000000101000111; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b01001011010111110000000000000101; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b00011111001100001001101000111100; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b01111110000101111010000111000011; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b00111000011101101010000110100101; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b00111001101000100100111011000010; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b01111000010011101110000110101000; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 6th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b10011001101101010000001100010000; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b10101001110001101001111111101010; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b11100000100100011110111110011010; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b10100100011100100110011101010000; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b11011110111000011111000010101101; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b10111000100110000111101001101100; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b11111110110010001100100111100100; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b01000000110011111011101110011101; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b00001011010010000110101001010100; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b01110001011001100011010110010100; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 7th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b11010111011110110110001110000111; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b00001101000101101010100001011011; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b11000010010100010000100000100000; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b00111111110100101010010101100111; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b10101011101111010000001101010001; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b00100101000000111011001000111101; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b10001010010001011111011100110011; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b10000001101001110010110100101000; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b01001111100110111011101110010010; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b11100101011110100101111011111001; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 8th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b00001101001111001000011010101010; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b00111010000001000010001111000011; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b10000110011010101100011100001110; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b10100101100111101111011011010110; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b10000111000111001100001111110001; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b10001001101100101100010011110100; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b10001110101010000100110100001100; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b10100000110101001011011011011110; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b01100001000000111010010001011000; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b10000110111001111010110100111111; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 9th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b11011111000010001100011001000100; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b00100100010001001001001011000101; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b01110011101101010000101101001010; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b01001110101110001000111111110011; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b10111000010101001001001010010000; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b10000010011001010010110001100111; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b10010011000010011110110010101000; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b10000111001101001011101100101111; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b00111110110010100001110101010001; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b11000100011011111101101001101100; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 10th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b11111010101001111111101001010000; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b01011011111000111110101010010000; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b10111000011001111100010110110011; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b10001101001100111101001011101110; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b00101100000110101101000010010110; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b00100011011101011010110011111111; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b10010001101001011011010101011111; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b10100000001001100011000111100011; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b01101010100111110100001110111001; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b01011010100101000000111111000011; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 11th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b11001101000000100101010001101100; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b11000010111000010011011010000000; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b11000011110110000110110000010111; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b11101101101010001010100101000011; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b11010011101110100010010110010001; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b10100110001111110110001000110111; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b10011000011001110111011000011100; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b01000101101100000001101100011101; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b01000000110001111010001010011110; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b01110111011111010101010000100101; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 12th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b01010101111011011100101000111111; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b10010011111001101101101011111001; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b11101000010001001010100110001101; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b01001000001111100101110010110101; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b10100011001100110100110101001101; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b01101001000111101100011000110000; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b11000011101010001111000100110010; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b00000001100111111101101100010000; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b11100001100001011101010101101000; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b11010100101111100000001001111110; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 13th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b00110011010000111111001110000001; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b01111100010010001010100100110011; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b11010100010110110100001100000001; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b11001110100001000111100111000011; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b00101110011100101100010110000011; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b01011000001111010100101100001101; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b00110001001011010011010111000100; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b00001001010010101110110101100000; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b11100110110010101011001011001011; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b10001001111111010101001001011101; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 14th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b00110001111111001000100011101100; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b00001110101110011000011010010010; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b00101000111011110000011111111101; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b01001111100110011110110011000011; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b00101000100011110001011100000011; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b01110011111111000000111001011001; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b01101001011010000111111111100100; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b00001100100001100011100110100011; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b10001011110000001010010101111111; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b00000111001110111001101011010010; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 15th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b11011011011001010010010100010001; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b00011000100111111110101011010100; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b01011100101111000010100100010010; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b01100110000111000100110100011100; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b10110111000100101111011110110010; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b10011011110110111100100010110101; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b11101010101011001000100000001011; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b10100111111010000011010000001010; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b10101110011000100111101110001001; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b11000110111010001101010001101100; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 16th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b11000110010101000100000000100100; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b10001101111110111100101010110001; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b01000000110110001000100001110110; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b11100000000000010111010101001100; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b01100111001000111001110110001001; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b00101101001110110110001111000010; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b00111000110111100111010000010011; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b10111110101010010001011110111001; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b10100010111111101011010010101001; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b01000110100000110100111010110100; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 17th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b10000100110100110101100111010100; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b00111010110001111010011010100001; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b01011011010101011111010101000011; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b11001101001011110111110111001101; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b11001111110111000010000011011101; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b00110011111110110110111111100111; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b00011100010011010110110001010101; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b10000110101000011111010101110100; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b11110011100000110101101111001101; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b01010011100111110101000100110011; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 18th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b10110100011000111101011001011010; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b00111100001011011111000100011110; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b00111010110100011110100000101101; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b01111011111001000011010101101010; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b10110100000001101011000001110001; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b00011100111010001001100101101011; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b01110001100100001010101010011001; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b01000000010101001101110100000101; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b01110011101001011100011011101001; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b00110101100001000000000001000001; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 19th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b10110100011111110100111001001111; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b11001000001001101111110101100001; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b01001110101111101101011101011110; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b10000101011101110110001000111001; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b00111100101001110111111001011000; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b10100000110001011000011000010011; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b01100100010101110010110100110001; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b11010100001111111111001000001011; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b10101100010110100010101101001010; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b11000110010001111010110001011111; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // 20th round:
            #36000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1280; ram_i_data1 = 32'b10001000111101000100000111101111; // action  31 ~   0
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1281; ram_i_data1 = 32'b11110010100000000110100001010100; // action  63 ~  32
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1282; ram_i_data1 = 32'b00010101100111001100001111001001; // action  95 ~  64
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1283; ram_i_data1 = 32'b10110100010011110001001001001000; // action 127 ~  96
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1284; ram_i_data1 = 32'b11000110011111001010001111011000; // action 159 ~ 128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1285; ram_i_data1 = 32'b10111000000100111011001011001000; // action 191 ~ 160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1286; ram_i_data1 = 32'b10100101011111001001010010100010; // action 223 ~ 192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1287; ram_i_data1 = 32'b11011010001101110111011011110000; // action 255 ~ 224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1288; ram_i_data1 = 32'b00000010100110100110010110100000; // action 287 ~ 256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1289; ram_i_data1 = 32'b10100111110110000001111000101001; // action 319 ~ 288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1290; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
    end

    // record observations
        integer fpga_ans;
        localparam FPGA_ANS_WD_NUM = SW_ENV_NUM*(u_Pipeline.DST_ENV_WD_NUM-2) +
                                    SW_ENV_NUM*u_Pipeline.RWD_WL/DATA_WL +
                                    SW_ENV_NUM/DATA_WL;
        initial begin
            fpga_ans = $fopen("/data0/FPGA_GYM/verilog/LocalStoreTemplate/LocalStoreTemplate.srcs/sim_1/new/fpga_ans.txt", "w");
            #640000 $fclose(fpga_ans);
        end
        always @(posedge new_round or negedge rstn) begin
            if (~rstn) begin
                cycle_cnt <= `ALL1(64);
            end else begin: write_fpga_ans
                reg [DATA_WL : 0] i;
                cycle_cnt <= cycle_cnt + 1;
                if (cycle_cnt[63] == 0) begin // there has been some result in BRAM
                    $fwrite(fpga_ans, "Iteration %d:\n", cycle_cnt);
                    for (i = `ZERO($clog2(SW_ENV_NUM)+1); i < FPGA_ANS_WD_NUM; i = i + 1) begin
                        $fwrite(fpga_ans, "%h%h%h%h ",
                                        u_My_RAM.Memory[u_Pipeline.OUT_INIT_ADDR+i][ 7: 0],
                                        u_My_RAM.Memory[u_Pipeline.OUT_INIT_ADDR+i][15: 8],
                                        u_My_RAM.Memory[u_Pipeline.OUT_INIT_ADDR+i][23:16],
                                        u_My_RAM.Memory[u_Pipeline.OUT_INIT_ADDR+i][31:24]);
                    end
                    $fwrite(fpga_ans, "\n\n");
                end
            end
        end

    // connect ports
        // cliffwalking_step inputs
            assign uut_i_data = ram_o_data2;
        // BRAM inputs
            assign ram_i_wr2   = ~&uut_o_wea;
            assign ram_i_addr2 = uut_o_addr[ADDR_WL-1:2];
            assign ram_i_data2 = uut_o_data;

    Pipeline #(.DATA_WL(DATA_WL), .ADDR_WL(ADDR_WL), .WEA_WL(WEA_WL), .SW_ENV_NUM(SW_ENV_NUM)) u_Pipeline(
        .i_clk  ( clk  ),
        .i_rstn ( rstn ),
        .i_data ( uut_i_data[DATA_WL-1:0] ),
        .o_data ( uut_o_data[DATA_WL-1:0] ),
        .o_addr ( uut_o_addr[ADDR_WL-1:0] ),
        .o_en   ( uut_o_en ),
        .o_wea  ( uut_o_wea[WEA_WL-1:0] ),
        .o_rstb ( uut_o_rstb )
    );
    My_RAM #(.ADDR_WIDTH(RAM_ADDR_WL), .DATA_WIDTH(DATA_WL)) u_My_RAM(
        .i_clk   ( clk ),
        .i_rstn  ( rstn ),
        .i_wr1   ( ram_i_wr1 ),
        .i_addr1 ( ram_i_addr1[RAM_ADDR_WL-1:0] ),
        .i_data1 ( ram_i_data1[DATA_WL-1:0] ),
        .o_data1 ( ram_o_data1[DATA_WL-1:0] ),
        .i_wr2   ( ram_i_wr2 ),
        .i_addr2 ( ram_i_addr2[RAM_ADDR_WL-1:0] ),
        .i_data2 ( ram_i_data2[DATA_WL-1:0] ),
        .o_data2 ( ram_o_data2[DATA_WL-1:0] )
    );

endmodule