`timescale 1ns / 1ps
`ifndef ONE // 1
`define ONE(WL) {{(WL-1){1'b0}}, 1'b1}
`endif

`ifndef ZERO // 0
`define ZERO(WL) {(WL){1'b0}}
`endif

`ifndef ALL1 // 111111
`define ALL1(WL) {(WL){1'b1}}
`endif

module Pipline_tb();

    parameter DATA_WL     = 32'd32;
    parameter ADDR_WL     = 32'd32;
    parameter WEA_WL      = 32'd4;
    parameter SW_ENV_NUM  = 30'd192;
    parameter RAM_ADDR_WL = 11; // if RAM_ADDR_WL is 32, simulation will be very slow 

    reg        clk = 0;
    reg        rstn;
    reg [63:0] clk_cnt;
    reg [63:0] cycle_cnt;

    reg new_round; // a new round of compute is started

    // Pipeline ports
        wire [DATA_WL-1:0] uut_i_data;
        wire [DATA_WL-1:0] uut_o_data;
        wire [ADDR_WL-1:0] uut_o_addr;
        wire               uut_o_en;
        wire [WEA_WL-1:0]  uut_o_wea;
        wire               uut_o_rstb;

    // BRAM ports
        reg                    ram_i_wr1;
        reg  [RAM_ADDR_WL-1:0] ram_i_addr1;
        reg  [DATA_WL-1:0]     ram_i_data1;
        wire [DATA_WL-1:0]     ram_o_data1;
        wire                   ram_i_wr2;
        wire [RAM_ADDR_WL-1:0] ram_i_addr2;
        wire [DATA_WL-1:0]     ram_i_data2;
        wire [DATA_WL-1:0]     ram_o_data2;

    always #5 clk = !clk;

    initial begin
        rstn = 1;
        #10 rstn = 0;
        #10 rstn = 1;
        // #10000 $finish;
    end

    always @(posedge clk or negedge rstn) begin
        if (rstn == 1'b0) begin
            clk_cnt <= 64'b0;
        end else begin
            clk_cnt <= clk_cnt + 1'b1;
        end
    end
    parameter MULTI_CLR = 0;
    generate
        if (MULTI_CLR == 1) begin
            initial begin // write initial data
                #0  ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0; ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 0:
                    // ENV   0:
                    #20 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 1:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 2:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 3:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 4:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 5:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 6:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 7:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 8:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 9:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 10:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 11:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 12:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 13:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 14:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 15:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 16:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 17:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 18:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 19:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 20:
                    // ENV   0:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
            end
        end else begin
            initial begin // write initial data
                #0  ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0; ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 0:
                    // ENV   0:
                    #20 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'h00000000;

                    // ENV   1:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'h00000000;

                    // ENV   2:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'h00000000;

                    // ENV   3:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h00000000;

                    // ENV   4:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h00000000;

                    // ENV   5:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'h00000000;

                    // ENV   6:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h00000000;

                    // ENV   7:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h00000000;

                    // ENV   8:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'h00000000;

                    // ENV   9:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'h00000000;

                    // ENV  10:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'h00000000;

                    // ENV  11:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h00000000;

                    // ENV  12:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h00000000;

                    // ENV  13:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h00000000;

                    // ENV  14:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h00000000;

                    // ENV  15:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h00000000;

                    // ENV  16:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'h00000000;

                    // ENV  17:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h00000000;

                    // ENV  18:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'h00000000;

                    // ENV  19:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'h00000000;

                    // ENV  20:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h00000000;

                    // ENV  21:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'h00000000;

                    // ENV  22:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'h00000000;

                    // ENV  23:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h00000000;

                    // ENV  24:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'h00000000;

                    // ENV  25:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'h00000000;

                    // ENV  26:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'h00000000;

                    // ENV  27:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h00000000;

                    // ENV  28:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'h00000000;

                    // ENV  29:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'h00000000;

                    // ENV  30:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h00000000;

                    // ENV  31:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h00000000;

                    // ENV  32:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h00000000;

                    // ENV  33:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'h00000000;

                    // ENV  34:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h00000000;

                    // ENV  35:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h00000000;

                    // ENV  36:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'h00000000;

                    // ENV  37:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'h00000000;

                    // ENV  38:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'h00000000;

                    // ENV  39:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h00000000;

                    // ENV  40:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h00000000;

                    // ENV  41:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'h00000000;

                    // ENV  42:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h00000000;

                    // ENV  43:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h00000000;

                    // ENV  44:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h00000000;

                    // ENV  45:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'h00000000;

                    // ENV  46:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'h00000000;

                    // ENV  47:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'h00000000;

                    // ENV  48:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h00000000;

                    // ENV  49:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'h00000000;

                    // ENV  50:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'h00000000;

                    // ENV  51:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'h00000000;

                    // ENV  52:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h00000000;

                    // ENV  53:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'h00000000;

                    // ENV  54:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h00000000;

                    // ENV  55:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h00000000;

                    // ENV  56:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h00000000;

                    // ENV  57:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'h00000000;

                    // ENV  58:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'h00000000;

                    // ENV  59:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h00000000;

                    // ENV  60:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h00000000;

                    // ENV  61:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h00000000;

                    // ENV  62:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'h00000000;

                    // ENV  63:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'h00000000;

                    // ENV  64:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h00000000;

                    // ENV  65:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h00000000;

                    // ENV  66:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'h00000000;

                    // ENV  67:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h00000000;

                    // ENV  68:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h00000000;

                    // ENV  69:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h00000000;

                    // ENV  70:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h00000000;

                    // ENV  71:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h00000000;

                    // ENV  72:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'h00000000;

                    // ENV  73:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'h00000000;

                    // ENV  74:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'h00000000;

                    // ENV  75:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h00000000;

                    // ENV  76:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h00000000;

                    // ENV  77:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h00000000;

                    // ENV  78:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h00000000;

                    // ENV  79:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h00000000;

                    // ENV  80:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h00000000;

                    // ENV  81:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h00000000;

                    // ENV  82:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h00000000;

                    // ENV  83:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h00000000;

                    // ENV  84:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h00000000;

                    // ENV  85:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h00000000;

                    // ENV  86:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h00000000;

                    // ENV  87:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h00000000;

                    // ENV  88:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h00000000;

                    // ENV  89:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h00000000;

                    // ENV  90:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h00000000;

                    // ENV  91:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h00000000;

                    // ENV  92:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h00000000;

                    // ENV  93:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h00000000;

                    // ENV  94:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h00000000;

                    // ENV  95:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h00000000;

                    // ENV  96:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h00000000;

                    // ENV  97:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h00000000;

                    // ENV  98:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h00000000;

                    // ENV  99:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h00000000;

                    // ENV 100:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h00000000;

                    // ENV 101:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h00000000;

                    // ENV 102:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h00000000;

                    // ENV 103:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h00000000;

                    // ENV 104:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h00000000;

                    // ENV 105:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h00000000;

                    // ENV 106:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h00000000;

                    // ENV 107:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h00000000;

                    // ENV 108:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h00000000;

                    // ENV 109:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h00000000;

                    // ENV 110:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h00000000;

                    // ENV 111:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h00000000;

                    // ENV 112:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h00000000;

                    // ENV 113:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h00000000;

                    // ENV 114:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h00000000;

                    // ENV 115:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd577; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd578; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd579; ram_i_data1 = 32'h00000000;

                    // ENV 116:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd580; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd581; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd582; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd583; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd584; ram_i_data1 = 32'h00000000;

                    // ENV 117:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd585; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd586; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd587; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd588; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd589; ram_i_data1 = 32'h00000000;

                    // ENV 118:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd590; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd591; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd592; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd593; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd594; ram_i_data1 = 32'h00000000;

                    // ENV 119:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd595; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd596; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd597; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd598; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd599; ram_i_data1 = 32'h00000000;

                    // ENV 120:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd600; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd601; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd602; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd603; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd604; ram_i_data1 = 32'h00000000;

                    // ENV 121:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd605; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd606; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd607; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd608; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd609; ram_i_data1 = 32'h00000000;

                    // ENV 122:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd610; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd611; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd612; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd613; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd614; ram_i_data1 = 32'h00000000;

                    // ENV 123:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd615; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd616; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd617; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd618; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd619; ram_i_data1 = 32'h00000000;

                    // ENV 124:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd620; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd621; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd622; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd623; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd624; ram_i_data1 = 32'h00000000;

                    // ENV 125:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd625; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd626; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd627; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd628; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd629; ram_i_data1 = 32'h00000000;

                    // ENV 126:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd630; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd631; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd632; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd633; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd634; ram_i_data1 = 32'h00000000;

                    // ENV 127:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd635; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd636; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd637; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd638; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd639; ram_i_data1 = 32'h00000000;

                    // ENV 128:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd640; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd641; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd642; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd643; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd644; ram_i_data1 = 32'h00000000;

                    // ENV 129:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd645; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd646; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd647; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd648; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd649; ram_i_data1 = 32'h00000000;

                    // ENV 130:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd650; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd651; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd652; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd653; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd654; ram_i_data1 = 32'h00000000;

                    // ENV 131:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd655; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd656; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd657; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd658; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd659; ram_i_data1 = 32'h00000000;

                    // ENV 132:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd660; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd661; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd662; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd663; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd664; ram_i_data1 = 32'h00000000;

                    // ENV 133:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd665; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd666; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd667; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd668; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd669; ram_i_data1 = 32'h00000000;

                    // ENV 134:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd670; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd671; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd672; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd673; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd674; ram_i_data1 = 32'h00000000;

                    // ENV 135:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd675; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd676; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd677; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd678; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd679; ram_i_data1 = 32'h00000000;

                    // ENV 136:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd680; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd681; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd682; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd683; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd684; ram_i_data1 = 32'h00000000;

                    // ENV 137:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd685; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd686; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd687; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd688; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd689; ram_i_data1 = 32'h00000000;

                    // ENV 138:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd690; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd691; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd692; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd693; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd694; ram_i_data1 = 32'h00000000;

                    // ENV 139:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd695; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd696; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd697; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd698; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd699; ram_i_data1 = 32'h00000000;

                    // ENV 140:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd700; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd701; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd702; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd703; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd704; ram_i_data1 = 32'h00000000;

                    // ENV 141:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd705; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd706; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd707; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd708; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd709; ram_i_data1 = 32'h00000000;

                    // ENV 142:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd710; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd711; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd712; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd713; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd714; ram_i_data1 = 32'h00000000;

                    // ENV 143:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd715; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd716; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd717; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd718; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd719; ram_i_data1 = 32'h00000000;

                    // ENV 144:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd720; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd721; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd722; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd723; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd724; ram_i_data1 = 32'h00000000;

                    // ENV 145:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd725; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd726; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd727; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd728; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd729; ram_i_data1 = 32'h00000000;

                    // ENV 146:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd730; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd731; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd732; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd733; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd734; ram_i_data1 = 32'h00000000;

                    // ENV 147:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd735; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd736; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd737; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd738; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd739; ram_i_data1 = 32'h00000000;

                    // ENV 148:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd740; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd741; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd742; ram_i_data1 = 32'h00700000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd743; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd744; ram_i_data1 = 32'h00000000;

                    // ENV 149:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd745; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd746; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd747; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd748; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd749; ram_i_data1 = 32'h00000000;

                    // ENV 150:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd750; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd751; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd752; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd753; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd754; ram_i_data1 = 32'h00000000;

                    // ENV 151:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd755; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd756; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd757; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd758; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd759; ram_i_data1 = 32'h00000000;

                    // ENV 152:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd760; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd761; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd762; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd763; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd764; ram_i_data1 = 32'h00000000;

                    // ENV 153:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd765; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd766; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd767; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd768; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd769; ram_i_data1 = 32'h00000000;

                    // ENV 154:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd770; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd771; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd772; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd773; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd774; ram_i_data1 = 32'h00000000;

                    // ENV 155:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd775; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd776; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd777; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd778; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd779; ram_i_data1 = 32'h00000000;

                    // ENV 156:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd780; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd781; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd782; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd783; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd784; ram_i_data1 = 32'h00000000;

                    // ENV 157:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd785; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd786; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd787; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd788; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd789; ram_i_data1 = 32'h00000000;

                    // ENV 158:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd790; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd791; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd792; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd793; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd794; ram_i_data1 = 32'h00000000;

                    // ENV 159:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd795; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd796; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd797; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd798; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd799; ram_i_data1 = 32'h00000000;

                    // ENV 160:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd800; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd801; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd802; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd803; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd804; ram_i_data1 = 32'h00000000;

                    // ENV 161:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd805; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd806; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd807; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd808; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd809; ram_i_data1 = 32'h00000000;

                    // ENV 162:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd810; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd811; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd812; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd813; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd814; ram_i_data1 = 32'h00000000;

                    // ENV 163:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd815; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd816; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd817; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd818; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd819; ram_i_data1 = 32'h00000000;

                    // ENV 164:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd820; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd821; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd822; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd823; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd824; ram_i_data1 = 32'h00000000;

                    // ENV 165:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd825; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd826; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd827; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd828; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd829; ram_i_data1 = 32'h00000000;

                    // ENV 166:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd830; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd831; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd832; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd833; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd834; ram_i_data1 = 32'h00000000;

                    // ENV 167:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd835; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd836; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd837; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd838; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd839; ram_i_data1 = 32'h00000000;

                    // ENV 168:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd840; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd841; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd842; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd843; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd844; ram_i_data1 = 32'h00000000;

                    // ENV 169:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd845; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd846; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd847; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd848; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd849; ram_i_data1 = 32'h00000000;

                    // ENV 170:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd850; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd851; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd852; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd853; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd854; ram_i_data1 = 32'h00000000;

                    // ENV 171:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd855; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd856; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd857; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd858; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd859; ram_i_data1 = 32'h00000000;

                    // ENV 172:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd860; ram_i_data1 = 32'h00000005;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd861; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd862; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd863; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd864; ram_i_data1 = 32'h00000000;

                    // ENV 173:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd865; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd866; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd867; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd868; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd869; ram_i_data1 = 32'h00000000;

                    // ENV 174:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd870; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd871; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd872; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd873; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd874; ram_i_data1 = 32'h00000000;

                    // ENV 175:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd875; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd876; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd877; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd878; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd879; ram_i_data1 = 32'h00000000;

                    // ENV 176:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd880; ram_i_data1 = 32'h00000009;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd881; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd882; ram_i_data1 = 32'h00a00000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd883; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd884; ram_i_data1 = 32'h00000000;

                    // ENV 177:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd885; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd886; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd887; ram_i_data1 = 32'h00800000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd888; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd889; ram_i_data1 = 32'h00000000;

                    // ENV 178:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd890; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd891; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd892; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd893; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd894; ram_i_data1 = 32'h00000000;

                    // ENV 179:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd895; ram_i_data1 = 32'h00000007;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd896; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd897; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd898; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd899; ram_i_data1 = 32'h00000000;

                    // ENV 180:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd900; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd901; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd902; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd903; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd904; ram_i_data1 = 32'h00000000;

                    // ENV 181:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd905; ram_i_data1 = 32'h00000008;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd906; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd907; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd908; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd909; ram_i_data1 = 32'h00000000;

                    // ENV 182:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd910; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd911; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd912; ram_i_data1 = 32'h00600000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd913; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd914; ram_i_data1 = 32'h00000000;

                    // ENV 183:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd915; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd916; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd917; ram_i_data1 = 32'h00900000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd918; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd919; ram_i_data1 = 32'h00000000;

                    // ENV 184:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd920; ram_i_data1 = 32'h00000004;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd921; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd922; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd923; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd924; ram_i_data1 = 32'h00000000;

                    // ENV 185:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd925; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd926; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd927; ram_i_data1 = 32'h00200000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd928; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd929; ram_i_data1 = 32'h00000000;

                    // ENV 186:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd930; ram_i_data1 = 32'h00000006;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd931; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd932; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd933; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd934; ram_i_data1 = 32'h00000000;

                    // ENV 187:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd935; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd936; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd937; ram_i_data1 = 32'h00100000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd938; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd939; ram_i_data1 = 32'h00000000;

                    // ENV 188:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd940; ram_i_data1 = 32'h00000001;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd941; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd942; ram_i_data1 = 32'h00400000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd943; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd944; ram_i_data1 = 32'h00000000;

                    // ENV 189:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd945; ram_i_data1 = 32'h0000000a;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd946; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd947; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd948; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd949; ram_i_data1 = 32'h00000000;

                    // ENV 190:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd950; ram_i_data1 = 32'h00000003;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd951; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd952; ram_i_data1 = 32'h00500000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd953; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd954; ram_i_data1 = 32'h00000000;

                    // ENV 191:
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd955; ram_i_data1 = 32'h00000002;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd956; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd957; ram_i_data1 = 32'h00300000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd958; ram_i_data1 = 32'h00000000;
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd959; ram_i_data1 = 32'h00000000;

                    #18 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01101100001110101011110000101101; // action  31 ~   0 ( 9.0299535e26)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001100100001010100011100101; // action  63 ~  32 (-6.424183e-14)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101011001001001001101010010100; // action  95 ~  64 ( 5.847902e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100111100100100000110010011001; // action 127 ~  96 ( 1.3793958e24)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011011100001100100010111000; // action 159 ~ 128 (-8.554368e-13)
                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011010010100101100000001111011; // action 191 ~ 160 ( 1.4830345e16)

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 1:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b10011111100000011011111000000001; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b11100001000110000000000100110000; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00011010110010110001100000011100; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b10011110010100000000101101001000; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b00111101101011011100010101010101; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b10011100111000001001000111110101; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 2:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b10011110001000100000011010100001; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10110000010011001100100011011001; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00011011111000110110010101110101; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b00110111011110000001111011010111; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b01001000011010001001011011000100; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b10111111110111000101110011101101; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 3:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01010110011100001010111000101011; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101101101100101101101100110001; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b10111010000011001000101010100010; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b00100011011100110111101001010011; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b00101110011011001010011011011001; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b00011111101110011010011011100011; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 4:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b00011011000111001010100111111111; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b11101101001101000010001101110001; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b10100100100010010000110011101110; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b00011100011111011000000101000111; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b01001011010111110000000000000101; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b00011111001100001001101000111100; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 5:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b10011001101101010000001100010000; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10101001110001101001111111101010; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b11100000100100011110111110011010; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b10100100011100100110011101010000; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b11011110111000011111000010101101; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b10111000100110000111101001101100; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 6:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b11010111011110110110001110000111; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b00001101000101101010100001011011; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b11000010010100010000100000100000; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b00111111110100101010010101100111; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10101011101111010000001101010001; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b00100101000000111011001000111101; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 7:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b00001101001111001000011010101010; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b00111010000001000010001111000011; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b10000110011010101100011100001110; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b10100101100111101111011011010110; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10000111000111001100001111110001; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b10001001101100101100010011110100; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 8:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b11011111000010001100011001000100; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b00100100010001001001001011000101; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b01110011101101010000101101001010; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01001110101110001000111111110011; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10111000010101001001001010010000; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b10000010011001010010110001100111; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 9:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b11111010101001111111101001010000; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b01011011111000111110101010010000; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b10111000011001111100010110110011; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b10001101001100111101001011101110; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b00101100000110101101000010010110; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b00100011011101011010110011111111; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 10:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b11001101000000100101010001101100; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b11000010111000010011011010000000; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b11000011110110000110110000010111; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b11101101101010001010100101000011; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b11010011101110100010010110010001; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b10100110001111110110001000110111; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 11:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b01010101111011011100101000111111; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10010011111001101101101011111001; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b11101000010001001010100110001101; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01001000001111100101110010110101; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10100011001100110100110101001101; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01101001000111101100011000110000; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 12:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b00110011010000111111001110000001; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b01111100010010001010100100110011; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b11010100010110110100001100000001; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b11001110100001000111100111000011; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b00101110011100101100010110000011; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01011000001111010100101100001101; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 13:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b00110001111111001000100011101100; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b00001110101110011000011010010010; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00101000111011110000011111111101; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01001111100110011110110011000011; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b00101000100011110001011100000011; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b01110011111111000000111001011001; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 14:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b11011011011001010010010100010001; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b00011000100111111110101011010100; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b01011100101111000010100100010010; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01100110000111000100110100011100; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10110111000100101111011110110010; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b10011011110110111100100010110101; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 15:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b11000110010101000100000000100100; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b10001101111110111100101010110001; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b01000000110110001000100001110110; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b11100000000000010111010101001100; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b01100111001000111001110110001001; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b00101101001110110110001111000010; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 16:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b10000100110100110101100111010100; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b00111010110001111010011010100001; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b01011011010101011111010101000011; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b11001101001011110111110111001101; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b11001111110111000010000011011101; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b00110011111110110110111111100111; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 17:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b10110100011000111101011001011010; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b00111100001011011111000100011110; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00111010110100011110100000101101; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b01111011111001000011010101101010; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b10110100000001101011000001110001; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b00011100111010001001100101101011; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 18:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b10110100011111110100111001001111; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b11001000001001101111110101100001; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b01001110101111101101011101011110; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b10000101011101110110001000111001; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b00111100101001110111111001011000; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b10100000110001011000011000010011; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
                // round 19:
                    #18000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd960; ram_i_data1 = 32'b10001000111101000100000111101111; // action  31 ~   0
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd961; ram_i_data1 = 32'b11110010100000000110100001010100; // action  63 ~  32
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd962; ram_i_data1 = 32'b00010101100111001100001111001001; // action  95 ~  64
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd963; ram_i_data1 = 32'b10110100010011110001001001001000; // action 127 ~  96
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd964; ram_i_data1 = 32'b11000110011111001010001111011000; // action 159 ~ 128
                    #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd965; ram_i_data1 = 32'b10111000000100111011001011001000; // action 191 ~ 160

                    #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd966; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
                    #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
            end
        end
    endgenerate

    // record observations
        integer fpga_ans;
        localparam RWD_WL = 2, ACT_WL = 1;
        localparam STA_WL = 160; // a multiple of DATA_WL
        localparam OBS_WL = 32;  // a multiple of DATA_WL
        localparam ENV_NUM = 32; // a multiple of DATA_WL and PE_NUM

        localparam SRC_ENV_WD_NUM  = 30'd6; // STA_WL/DATA_WL + 1
        localparam DST_ENV_WD_NUM  = 30'd3; // OBS_WL/DATA_WL + 2
        localparam ACT_INIT_ADDR   = SW_ENV_NUM*(SRC_ENV_WD_NUM-1);
        localparam START_FLAG_ADDR = ACT_INIT_ADDR + (SW_ENV_NUM*ACT_WL/DATA_WL);
        localparam OUT_INIT_ADDR   = START_FLAG_ADDR + 1;
        localparam RWD_INIT_ADDR   = SW_ENV_NUM*(DST_ENV_WD_NUM-2);
        localparam DONE_INIT_ADDR  = RWD_INIT_ADDR + SW_ENV_NUM*RWD_WL/DATA_WL;
        localparam FPGA_ANS_WD_NUM = SW_ENV_NUM*(DST_ENV_WD_NUM-2) +
                                     SW_ENV_NUM*RWD_WL/DATA_WL +
                                     SW_ENV_NUM/DATA_WL;
        initial begin
            fpga_ans = $fopen("/data0/FPGA_GYM/verilog/BlackJack/BlackJack.srcs/sim_1/new/fpga_ans.txt", "w");
            #640000 $fclose(fpga_ans);
        end
        always @(posedge new_round or negedge rstn) begin
            if (~rstn) begin
                cycle_cnt <= `ALL1(64);
            end else begin: write_fpga_ans
                reg [DATA_WL : 0] i;
                cycle_cnt <= cycle_cnt + 1;
                if (cycle_cnt[63] == 0) begin // there has been some result in BRAM
                    $fwrite(fpga_ans, "Iteration %d:\n", cycle_cnt);
                    for (i = `ZERO($clog2(SW_ENV_NUM)+1); i < FPGA_ANS_WD_NUM; i = i + 1) begin
                        $fwrite(fpga_ans, "%h%h%h%h ",
                                        u_My_RAM.Memory[OUT_INIT_ADDR+i][ 7: 0],
                                        u_My_RAM.Memory[OUT_INIT_ADDR+i][15: 8],
                                        u_My_RAM.Memory[OUT_INIT_ADDR+i][23:16],
                                        u_My_RAM.Memory[OUT_INIT_ADDR+i][31:24]);
                    end
                    $fwrite(fpga_ans, "\n\n");
                end
            end
        end

    // connect ports
        // cliffwalking_step inputs
            assign uut_i_data = ram_o_data2;
        // BRAM inputs
            assign ram_i_wr2   = ~&uut_o_wea;
            assign ram_i_addr2 = uut_o_addr[ADDR_WL-1:2];
            assign ram_i_data2 = uut_o_data;

    Pipeline #(.DATA_WL(DATA_WL), .ADDR_WL(ADDR_WL), .WEA_WL(WEA_WL), .SW_ENV_NUM(SW_ENV_NUM)) u_Pipeline(
        .i_clk  ( clk  ),
        .i_rstn ( rstn ),
        .i_data ( uut_i_data[DATA_WL-1:0] ),
        .o_data ( uut_o_data[DATA_WL-1:0] ),
        .o_addr ( uut_o_addr[ADDR_WL-1:0] ),
        .o_en   ( uut_o_en ),
        .o_wea  ( uut_o_wea[WEA_WL-1:0] ),
        .o_rstb ( uut_o_rstb ),
        .i_debug ( 13'b00000_00000100 ),
        .o_debug ()
    );
    My_RAM #(.ADDR_WIDTH(RAM_ADDR_WL), .DATA_WIDTH(DATA_WL)) u_My_RAM(
        .i_clk   ( clk ),
        .i_rstn  ( rstn ),
        .i_wr1   ( ram_i_wr1 ),
        .i_addr1 ( ram_i_addr1[RAM_ADDR_WL-1:0] ),
        .i_data1 ( ram_i_data1[DATA_WL-1:0] ),
        .o_data1 ( ram_o_data1[DATA_WL-1:0] ),
        .i_wr2   ( ram_i_wr2 ),
        .i_addr2 ( ram_i_addr2[RAM_ADDR_WL-1:0] ),
        .i_data2 ( ram_i_data2[DATA_WL-1:0] ),
        .o_data2 ( ram_o_data2[DATA_WL-1:0] )
    );

endmodule