`timescale 1ns / 1ps
`ifndef ONE // 1
`define ONE(WL) {{(WL-1){1'b0}}, 1'b1}
`endif

`ifndef ZERO // 0
`define ZERO(WL) {(WL){1'b0}}
`endif

`ifndef ALL1 // 111111
`define ALL1(WL) {(WL){1'b1}}
`endif

module Pipline_tb();

    parameter DATA_WL = 32'd32;
    parameter ADDR_WL = 32'd32;
    parameter WEA_WL  = 32'd4;
    parameter SW_ENV_NUM = 30'd192;
    parameter RAM_ADDR_WL = 12; // if RAM_ADDR_WL is 32, simulation will be very slow 

    reg        clk = 0;
    reg        rstn;
    reg [63:0] clk_cnt;
    reg [63:0] cycle_cnt;

    reg new_round; // a new round of compute is started

    // Pipeline ports
        wire [DATA_WL-1:0] uut_i_data;
        wire [DATA_WL-1:0] uut_o_data;
        wire [ADDR_WL-1:0] uut_o_addr;
        wire               uut_o_en;
        wire [WEA_WL-1:0]  uut_o_wea;
        wire               uut_o_rstb;

    // BRAM ports
        reg                    ram_i_wr1;
        reg  [RAM_ADDR_WL-1:0] ram_i_addr1;
        reg  [DATA_WL-1:0]     ram_i_data1;
        wire [DATA_WL-1:0]     ram_o_data1;
        wire                   ram_i_wr2;
        wire [RAM_ADDR_WL-1:0] ram_i_addr2;
        wire [DATA_WL-1:0]     ram_i_data2;
        wire [DATA_WL-1:0]     ram_o_data2;

    always #5 clk = !clk;

    initial begin
        rstn = 1;
        #10 rstn = 0;
        #10 rstn = 1;
    //  #10000 $finish;
    end

    always @(posedge clk or negedge rstn) begin
        if (rstn == 1'b0) begin
            clk_cnt <= 64'b0;
        end else begin
            clk_cnt <= clk_cnt + 1'b1;
        end
    end
    initial begin // write initial data
        #0  ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0; ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 0:
            #20 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd0; ram_i_data1 = 32'hbef42995; // θ0:-0.47687975
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd1; ram_i_data1 = 32'hbfdd3a26; // ω0:-1.72833705

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd2; ram_i_data1 = 32'h402e0ca8; // θ1: 2.71952248
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd3; ram_i_data1 = 32'hbf6305ee; // ω1:-0.88680923

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd4; ram_i_data1 = 32'hbf206b33; // θ2:-0.62663573
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd5; ram_i_data1 = 32'hbeaa2940; // ω2:-0.33234596

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd6; ram_i_data1 = 32'h3da1fa47; // θ3: 0.07909065
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd7; ram_i_data1 = 32'h3e1a25d1; // ω3: 0.15053488

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd8; ram_i_data1 = 32'h400e520d; // θ4: 2.22375798
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd9; ram_i_data1 = 32'hc023134c; // ω4:-2.54805279

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd10; ram_i_data1 = 32'h40043306; // θ5: 2.06561422
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd11; ram_i_data1 = 32'h40058199; // ω5: 2.08603501

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd12; ram_i_data1 = 32'h3f0910ae; // θ6: 0.53541076
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd13; ram_i_data1 = 32'hbd3cfc9b; // ω6:-0.04613934

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd14; ram_i_data1 = 32'hbf4646ca; // θ7:-0.77451766
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd15; ram_i_data1 = 32'h40253ee5; // ω7: 2.58196378

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd16; ram_i_data1 = 32'hbf56d2f3; // θ8:-0.83915633
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd17; ram_i_data1 = 32'h3fb751a8; // ω8: 1.43217945

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd18; ram_i_data1 = 32'h3e475d84; // θ9: 0.19469267
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd19; ram_i_data1 = 32'h3ffb2db7; // ω9: 1.96233261

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd20; ram_i_data1 = 32'hc01d7954; // θ10:-2.46053028
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd21; ram_i_data1 = 32'h400aeadf; // ω10: 2.17058539

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd22; ram_i_data1 = 32'h3fe89178; // θ11: 1.81693935
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd23; ram_i_data1 = 32'h3ea3db02; // ω11: 0.32003027

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd24; ram_i_data1 = 32'h3fd7bebd; // θ12: 1.68550837
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd25; ram_i_data1 = 32'hbf03c40f; // ω12:-0.51471037

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd26; ram_i_data1 = 32'h400cd37a; // θ13: 2.20040751
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd27; ram_i_data1 = 32'hc0161d4e; // ω13:-2.34553862

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd28; ram_i_data1 = 32'h3e147070; // θ14: 0.14496017
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd29; ram_i_data1 = 32'hc0341714; // ω14:-2.81390858

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd30; ram_i_data1 = 32'h4009630c; // θ15: 2.14667034
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd31; ram_i_data1 = 32'h3f82add6; // ω15: 1.02093005

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd32; ram_i_data1 = 32'hbff9fb2b; // θ16:-1.95297754
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd33; ram_i_data1 = 32'h3f651fa2; // ω16: 0.89501393

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd34; ram_i_data1 = 32'h40374ef8; // θ17: 2.86419487
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd35; ram_i_data1 = 32'hc02a11ae; // ω17:-2.65732908

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd36; ram_i_data1 = 32'hc01fd41b; // θ18:-2.49732089
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd37; ram_i_data1 = 32'hc01fb723; // ω18:-2.49555278

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd38; ram_i_data1 = 32'hbcd313b2; // θ19:-0.02576623
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd39; ram_i_data1 = 32'h4000ab2a; // ω19: 2.01044703

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd40; ram_i_data1 = 32'hbfa5b46b; // θ20:-1.29456842
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd41; ram_i_data1 = 32'h402e8494; // ω20: 2.72684193

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd42; ram_i_data1 = 32'h3ec7c722; // θ21: 0.39019114
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd43; ram_i_data1 = 32'hbea85d77; // ω21:-0.32883808

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd44; ram_i_data1 = 32'hbff0a1a7; // θ22:-1.87993324
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd45; ram_i_data1 = 32'h3a2f77b0; // ω22: 0.00066936

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd46; ram_i_data1 = 32'h4014ff42; // θ23: 2.32807970
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd47; ram_i_data1 = 32'hbf7d5abc; // ω23:-0.98966575

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd48; ram_i_data1 = 32'h3f6deb52; // θ24: 0.92937195
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd49; ram_i_data1 = 32'hc043198b; // ω24:-3.04843402

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd50; ram_i_data1 = 32'hbf6d5f29; // θ25:-0.92723328
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd51; ram_i_data1 = 32'h4000363e; // ω25: 2.00331068

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd52; ram_i_data1 = 32'hbf2c8239; // θ26:-0.67386204
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd53; ram_i_data1 = 32'h4046cc86; // ω26: 3.10623312

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd54; ram_i_data1 = 32'hc020a554; // θ27:-2.51009083
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd55; ram_i_data1 = 32'hbe4a7b8e; // ω27:-0.19773695

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd56; ram_i_data1 = 32'h3fb67793; // θ28: 1.42552412
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd57; ram_i_data1 = 32'h40324767; // ω28: 2.78560805

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd58; ram_i_data1 = 32'hc0191cfc; // θ29:-2.39239407
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd59; ram_i_data1 = 32'h400e99d6; // ω29: 2.22813940

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd60; ram_i_data1 = 32'hc0412a5b; // θ30:-3.01821017
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd61; ram_i_data1 = 32'hbe42cf1d; // ω30:-0.19024320

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd62; ram_i_data1 = 32'h3ef4a9a6; // θ31: 0.47785681
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd63; ram_i_data1 = 32'hbe38fea2; // ω31:-0.18065885

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd64; ram_i_data1 = 32'h3f8497d7; // θ32: 1.03588378
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd65; ram_i_data1 = 32'hbffb7c29; // ω32:-1.96472657

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd66; ram_i_data1 = 32'h3fe89fa7; // θ33: 1.81737220
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd67; ram_i_data1 = 32'hbf03b9c6; // ω33:-0.51455343

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd68; ram_i_data1 = 32'h3cb0a1a0; // θ34: 0.02156144
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd69; ram_i_data1 = 32'h3ff5244b; // ω34: 1.91517007

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd70; ram_i_data1 = 32'hc01c167e; // θ35:-2.43887281
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd71; ram_i_data1 = 32'h3f1a6087; // ω35: 0.60303539

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd72; ram_i_data1 = 32'h3f8eff43; // θ36: 1.11716497
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd73; ram_i_data1 = 32'h40119097; // ω36: 2.27445006

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd74; ram_i_data1 = 32'h403c1e90; // θ37: 2.93936539
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd75; ram_i_data1 = 32'hc006b85c; // ω37:-2.10500240

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd76; ram_i_data1 = 32'h3f3c68ec; // θ38: 0.73597598
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd77; ram_i_data1 = 32'hbfee0255; // ω38:-1.85944617

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd78; ram_i_data1 = 32'hbfed6516; // θ39:-1.85464740
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd79; ram_i_data1 = 32'h3ec4fd40; // ω39: 0.38474464

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd80; ram_i_data1 = 32'h400097cb; // θ40: 2.00926471
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd81; ram_i_data1 = 32'h4037192c; // ω40: 2.86091137

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd82; ram_i_data1 = 32'h4042c5bd; // θ41: 3.04331899
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd83; ram_i_data1 = 32'hbf91ccf2; // ω41:-1.13906693

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd84; ram_i_data1 = 32'hbfe77690; // θ42:-1.80830574
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd85; ram_i_data1 = 32'h3f7b4e33; // ω42: 0.98166198

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd86; ram_i_data1 = 32'hc0334959; // θ43:-2.80135179
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd87; ram_i_data1 = 32'hbd8fda9f; // ω43:-0.07024121

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd88; ram_i_data1 = 32'hbfbcf032; // θ44:-1.47608018
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd89; ram_i_data1 = 32'h3fde65c9; // ω44: 1.73748124

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd90; ram_i_data1 = 32'h3f78c318; // θ45: 0.97172689
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd91; ram_i_data1 = 32'h4007309c; // ω45: 2.11234188

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd92; ram_i_data1 = 32'hc02d5634; // θ46:-2.70838642
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd93; ram_i_data1 = 32'h3f764f88; // ω46: 0.96215105

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd94; ram_i_data1 = 32'hbe04643a; // θ47:-0.12928858
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd95; ram_i_data1 = 32'h40144363; // ω47: 2.31661296

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd96; ram_i_data1 = 32'h401f6123; // θ48: 2.49030375
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd97; ram_i_data1 = 32'hbe8a3b50; // ω48:-0.26998377

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd98; ram_i_data1 = 32'h3f9b0ccc; // θ49: 1.21132803
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd99; ram_i_data1 = 32'hbffd8e82; // ω49:-1.98091149

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd100; ram_i_data1 = 32'hbff45d2f; // θ50:-1.90909374
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd101; ram_i_data1 = 32'hbfc9488b; // ω50:-1.57252634

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd102; ram_i_data1 = 32'hc026d9a2; // θ51:-2.60703325
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd103; ram_i_data1 = 32'h3f74909c; // ω51: 0.95533156

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd104; ram_i_data1 = 32'h3f4a112a; // θ52: 0.78932440
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd105; ram_i_data1 = 32'hbfdfc483; // ω52:-1.74818456

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd106; ram_i_data1 = 32'hc00f31bb; // θ53:-2.23741031
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd107; ram_i_data1 = 32'hbfc34177; // ω53:-1.52543533

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd108; ram_i_data1 = 32'h3fc627c3; // θ54: 1.54808843
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd109; ram_i_data1 = 32'hc0342a6d; // ω54:-2.81508946

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd110; ram_i_data1 = 32'hbf97a7e7; // θ55:-1.18481147
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd111; ram_i_data1 = 32'hbf8e45ff; // ω55:-1.11151111

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd112; ram_i_data1 = 32'h40132eb6; // θ56: 2.29972601
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd113; ram_i_data1 = 32'hbfbe801e; // ω56:-1.48828483

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd114; ram_i_data1 = 32'hbf99206b; // θ57:-1.19630182
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd115; ram_i_data1 = 32'hc02bd2a2; // ω57:-2.68473101

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd116; ram_i_data1 = 32'h402bd5ac; // θ58: 2.68491650
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd117; ram_i_data1 = 32'hbe413d18; // ω58:-0.18870962

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd118; ram_i_data1 = 32'hbd579bae; // θ59:-0.05263870
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd119; ram_i_data1 = 32'h3fb478d2; // ω59: 1.40993714

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd120; ram_i_data1 = 32'h3ec00792; // θ60: 0.37505776
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd121; ram_i_data1 = 32'h401f70f8; // ω60: 2.49127007

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd122; ram_i_data1 = 32'h3fd19122; // θ61: 1.63724160
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd123; ram_i_data1 = 32'hc029a225; // ω61:-2.65052152

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd124; ram_i_data1 = 32'hbf5ff0f5; // θ62:-0.87477046
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd125; ram_i_data1 = 32'h3f461bec; // ω62: 0.77386355

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd126; ram_i_data1 = 32'hbff4cc29; // θ63:-1.91248047
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd127; ram_i_data1 = 32'hc012e87d; // ω63:-2.29543996

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd128; ram_i_data1 = 32'hbff267fc; // θ64:-1.89379835
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd129; ram_i_data1 = 32'hbf9da98e; // ω64:-1.23173690

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd130; ram_i_data1 = 32'hc02d4acf; // θ65:-2.70769095
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd131; ram_i_data1 = 32'hbff5feb0; // ω65:-1.92183495

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd132; ram_i_data1 = 32'hc00ceb5d; // θ66:-2.20186543
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd133; ram_i_data1 = 32'h3ff81b60; // ω66: 1.93833542

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd134; ram_i_data1 = 32'hc00a8d55; // θ67:-2.16487622
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd135; ram_i_data1 = 32'hbfdbd9f0; // ω67:-1.71758842

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd136; ram_i_data1 = 32'hbf8ae775; // θ68:-1.08518851
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd137; ram_i_data1 = 32'hbff1eb14; // ω68:-1.88998652

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd138; ram_i_data1 = 32'h3fb5f8cc; // θ69: 1.42165518
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd139; ram_i_data1 = 32'h3fc33302; // ω69: 1.52499413

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd140; ram_i_data1 = 32'h3e7443fd; // θ70: 0.23854060
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd141; ram_i_data1 = 32'hc03a0485; // ω70:-2.90652585

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd142; ram_i_data1 = 32'h3f740ed4; // θ71: 0.95335126
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd143; ram_i_data1 = 32'h3f65a1b8; // ω71: 0.89699888

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd144; ram_i_data1 = 32'hc02c876a; // θ72:-2.69576502
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd145; ram_i_data1 = 32'hbfd7f00f; // ω72:-1.68701351

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd146; ram_i_data1 = 32'h40464869; // θ73: 3.09816957
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd147; ram_i_data1 = 32'h3fb58a71; // ω73: 1.41828740

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd148; ram_i_data1 = 32'h3f5fddc1; // θ74: 0.87447745
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd149; ram_i_data1 = 32'hbde23a4e; // ω74:-0.11046277

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd150; ram_i_data1 = 32'hbf191fe4; // θ75:-0.59814286
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd151; ram_i_data1 = 32'hbe318099; // ω75:-0.17334212

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd152; ram_i_data1 = 32'hbf68a5e9; // θ76:-0.90878159
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd153; ram_i_data1 = 32'hbf3835bd; // ω76:-0.71956998

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd154; ram_i_data1 = 32'h3f21767f; // θ77: 0.63071436
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd155; ram_i_data1 = 32'h3f3f329c; // ω77: 0.74686599

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd156; ram_i_data1 = 32'hc0449cf6; // θ78:-3.07208014
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd157; ram_i_data1 = 32'hbea4f53d; // ω78:-0.32218352

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd158; ram_i_data1 = 32'hc00e95d4; // θ79:-2.22789478
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd159; ram_i_data1 = 32'h4033b915; // ω79: 2.80817151

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd160; ram_i_data1 = 32'h3e0f1468; // θ80: 0.13972628
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd161; ram_i_data1 = 32'hbfa569e6; // ω80:-1.29229426

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd162; ram_i_data1 = 32'hc04328c4; // θ81:-3.04936314
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd163; ram_i_data1 = 32'hbfd0d3bb; // ω81:-1.63146150

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd164; ram_i_data1 = 32'h3f8694db; // θ82: 1.05141771
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd165; ram_i_data1 = 32'h3fb8a926; // ω82: 1.44266200

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd166; ram_i_data1 = 32'hbe7c9dac; // θ83:-0.24669522
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd167; ram_i_data1 = 32'hc0056b89; // ω83:-2.08468843

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd168; ram_i_data1 = 32'h3fa7082b; // θ84: 1.30493677
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd169; ram_i_data1 = 32'hbfe59a57; // ω84:-1.79377258

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd170; ram_i_data1 = 32'h3f2de060; // θ85: 0.67920494
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd171; ram_i_data1 = 32'h3ef32332; // ω85: 0.47487789

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd172; ram_i_data1 = 32'h3fc7940a; // θ86: 1.55920529
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd173; ram_i_data1 = 32'h3f4b19a8; // ω86: 0.79336023

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd174; ram_i_data1 = 32'h3f14b53e; // θ87: 0.58089054
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd175; ram_i_data1 = 32'hc013ab7c; // ω87:-2.30734158

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd176; ram_i_data1 = 32'hc03f1521; // θ88:-2.98566461
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd177; ram_i_data1 = 32'h402b46b8; // ω88: 2.67619133

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd178; ram_i_data1 = 32'hbe247440; // θ89:-0.16059971
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd179; ram_i_data1 = 32'h40460ace; // ω89: 3.09440947

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd180; ram_i_data1 = 32'hbfd922dc; // θ90:-1.69637632
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd181; ram_i_data1 = 32'hbf4c0a75; // ω90:-0.79703456

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd182; ram_i_data1 = 32'hc03fcf24; // θ91:-2.99701786
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd183; ram_i_data1 = 32'hbf657d10; // ω91:-0.89643955

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd184; ram_i_data1 = 32'hc0341365; // θ92:-2.81368375
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd185; ram_i_data1 = 32'hbfc77598; // ω92:-1.55827618

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd186; ram_i_data1 = 32'hbefb45ef; // θ93:-0.49076793
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd187; ram_i_data1 = 32'hbfab504d; // ω93:-1.33838809

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd188; ram_i_data1 = 32'hc03d6720; // θ94:-2.95941925
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd189; ram_i_data1 = 32'hbf8bbca0; // ω94:-1.09169388

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd190; ram_i_data1 = 32'hbfc4668e; // θ95:-1.53437972
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd191; ram_i_data1 = 32'h3f30d4ba; // ω95: 0.69074595

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd192; ram_i_data1 = 32'hc0338e58; // θ96:-2.80556297
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd193; ram_i_data1 = 32'h40070e0b; // ω96: 2.11023211

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd194; ram_i_data1 = 32'hbfc3376a; // θ97:-1.52512860
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd195; ram_i_data1 = 32'hbe76baac; // ω97:-0.24094647

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd196; ram_i_data1 = 32'h3f365cdb; // θ98: 0.71235436
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd197; ram_i_data1 = 32'hbfe05cc1; // ω98:-1.75283062

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd198; ram_i_data1 = 32'h40090402; // θ99: 2.14086962
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd199; ram_i_data1 = 32'h3fe4c1d0; // ω99: 1.78716469

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd200; ram_i_data1 = 32'hbf8968ba; // θ100:-1.07350850
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd201; ram_i_data1 = 32'hc025e733; // ω100:-2.59223628

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd202; ram_i_data1 = 32'hbed27bb2; // θ101:-0.41109997
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd203; ram_i_data1 = 32'h3ef251b2; // ω101: 0.47327954

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd204; ram_i_data1 = 32'h4039dd88; // θ102: 2.90414619
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd205; ram_i_data1 = 32'hc00dd7f6; // ω102:-2.21630621

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd206; ram_i_data1 = 32'hbf810cb1; // θ103:-1.00819981
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd207; ram_i_data1 = 32'h3fe174a6; // ω103: 1.76137233

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd208; ram_i_data1 = 32'h3d6d5bb3; // θ104: 0.05794878
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd209; ram_i_data1 = 32'hbf0a7472; // ω104:-0.54083931

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd210; ram_i_data1 = 32'h4026e7b8; // θ105: 2.60789299
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd211; ram_i_data1 = 32'hbf863e11; // ω105:-1.04876912

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd212; ram_i_data1 = 32'hbf0c90b2; // θ106:-0.54908288
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd213; ram_i_data1 = 32'hc0376d2d; // ω106:-2.86603856

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd214; ram_i_data1 = 32'h3f9f4f7f; // θ107: 1.24461353
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd215; ram_i_data1 = 32'h3fcb2cee; // ω107: 1.58730865

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd216; ram_i_data1 = 32'hc014b3b6; // θ108:-2.32346869
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd217; ram_i_data1 = 32'h3fda90e2; // ω108: 1.70754647

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd218; ram_i_data1 = 32'h3ffccb43; // θ109: 1.97495306
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd219; ram_i_data1 = 32'h3f5eac21; // ω109: 0.86981398

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd220; ram_i_data1 = 32'h40454d6f; // θ110: 3.08285117
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd221; ram_i_data1 = 32'h3f48a0af; // ω110: 0.78370184

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd222; ram_i_data1 = 32'h3e885fe7; // θ111: 0.26635668
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd223; ram_i_data1 = 32'hbfafbb32; // ω111:-1.37290025

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd224; ram_i_data1 = 32'h3feba269; // θ112: 1.84089386
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd225; ram_i_data1 = 32'h400fb6c1; // ω112: 2.24552941

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd226; ram_i_data1 = 32'hbf9df878; // θ113:-1.23414516
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd227; ram_i_data1 = 32'h3faf9568; // ω113: 1.37174702

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd228; ram_i_data1 = 32'hc01dab0b; // θ114:-2.46356463
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd229; ram_i_data1 = 32'hbdd2dc58; // ω114:-0.10295933

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd230; ram_i_data1 = 32'hc038e06e; // θ115:-2.88869810
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd231; ram_i_data1 = 32'h403de278; // ω115: 2.96694756

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd232; ram_i_data1 = 32'hc013004c; // θ116:-2.29689312
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd233; ram_i_data1 = 32'h3f6da874; // ω116: 0.92835164

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd234; ram_i_data1 = 32'hbfecaa3e; // θ117:-1.84894538
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd235; ram_i_data1 = 32'h4029111b; // ω117: 2.64166903

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd236; ram_i_data1 = 32'hbfd0381f; // θ118:-1.62671268
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd237; ram_i_data1 = 32'hc000b281; // ω118:-2.01089501

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd238; ram_i_data1 = 32'hbfc2b544; // θ119:-1.52115679
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd239; ram_i_data1 = 32'hc042fdac; // ω119:-3.04673290

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd240; ram_i_data1 = 32'h3f8ad59e; // θ120: 1.08464408
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd241; ram_i_data1 = 32'h3f6cb1d5; // ω120: 0.92458850

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd242; ram_i_data1 = 32'h401bcbc9; // θ121: 2.43431306
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd243; ram_i_data1 = 32'h4009538f; // ω121: 2.14572501

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd244; ram_i_data1 = 32'h3f9c5fdd; // θ122: 1.22167552
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd245; ram_i_data1 = 32'h3f03d3cf; // ω122: 0.51495069

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd246; ram_i_data1 = 32'hbf84f422; // θ123:-1.03870034
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd247; ram_i_data1 = 32'h4016b002; // ω123: 2.35449266

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd248; ram_i_data1 = 32'hc0290278; // θ124:-2.64077568
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd249; ram_i_data1 = 32'hbf86cac9; // ω124:-1.05306351

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd250; ram_i_data1 = 32'hc03937f2; // θ125:-2.89403963
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd251; ram_i_data1 = 32'hbe982cf3; // ω125:-0.29721794

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd252; ram_i_data1 = 32'hbfefdf1e; // θ126:-1.87399650
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd253; ram_i_data1 = 32'h3e7b2d59; // ω126: 0.24529018

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd254; ram_i_data1 = 32'hbf26f75a; // θ127:-0.65221179
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd255; ram_i_data1 = 32'h40024ba6; // ω127: 2.03586721

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd256; ram_i_data1 = 32'h403930d1; // θ128: 2.89360452
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd257; ram_i_data1 = 32'hbfa06949; // ω128:-1.25321305

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd258; ram_i_data1 = 32'hbfc1c7f1; // θ129:-1.51391423
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd259; ram_i_data1 = 32'hbe3ba87c; // ω129:-0.18325990

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd260; ram_i_data1 = 32'h3f623d73; // θ130: 0.88375014
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd261; ram_i_data1 = 32'h40108f41; // ω130: 2.25874352

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd262; ram_i_data1 = 32'hc0185e33; // θ131:-2.38074946
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd263; ram_i_data1 = 32'hbfe02f95; // ω131:-1.75145209

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd264; ram_i_data1 = 32'h3eee75e3; // θ132: 0.46574315
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd265; ram_i_data1 = 32'h3fd28524; // ω132: 1.64468813

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd266; ram_i_data1 = 32'hbe3ac19a; // θ133:-0.18237916
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd267; ram_i_data1 = 32'h3f83d57e; // ω133: 1.02995276

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd268; ram_i_data1 = 32'h3eb20e8f; // θ134: 0.34776732
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd269; ram_i_data1 = 32'hbfcb871f; // ω134:-1.59006107

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd270; ram_i_data1 = 32'hc00e60fb; // θ135:-2.22466922
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd271; ram_i_data1 = 32'hbf542563; // ω135:-0.82869548

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd272; ram_i_data1 = 32'hc0135e2a; // θ136:-2.30262232
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd273; ram_i_data1 = 32'h402e290e; // ω136: 2.72125578

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd274; ram_i_data1 = 32'h4046706b; // θ137: 3.10061145
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd275; ram_i_data1 = 32'hc03ff9bb; // ω137:-2.99961734

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd276; ram_i_data1 = 32'h3cf1de61; // θ138: 0.02952498
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd277; ram_i_data1 = 32'hbffade58; // ω138:-1.95991039

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd278; ram_i_data1 = 32'hc048a78b; // θ139:-3.13522601
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd279; ram_i_data1 = 32'h3f7c485b; // ω139: 0.98547906

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd280; ram_i_data1 = 32'h40018aaa; // θ140: 2.02408838
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd281; ram_i_data1 = 32'hbfe45f73; // ω140:-1.78416288

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd282; ram_i_data1 = 32'h3d6abf79; // θ141: 0.05731151
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd283; ram_i_data1 = 32'hbf9363ca; // ω141:-1.15148282

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd284; ram_i_data1 = 32'h401dbdb1; // θ142: 2.46470284
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd285; ram_i_data1 = 32'hbfe5a7c9; // ω142:-1.79418290

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd286; ram_i_data1 = 32'hbf88244a; // θ143:-1.06360745
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd287; ram_i_data1 = 32'hc02ee7a5; // ω143:-2.73288846

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd288; ram_i_data1 = 32'h3f5e8e05; // θ144: 0.86935455
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd289; ram_i_data1 = 32'hbf8c9f51; // ω144:-1.09861195

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd290; ram_i_data1 = 32'h3fe2e964; // θ145: 1.77274752
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd291; ram_i_data1 = 32'h3f40e197; // ω145: 0.75344223

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd292; ram_i_data1 = 32'hbef5ffcf; // θ146:-0.48046729
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd293; ram_i_data1 = 32'hc0144561; // ω146:-2.31673455

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd294; ram_i_data1 = 32'hbf81bc7c; // θ147:-1.01356459
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd295; ram_i_data1 = 32'h3fb111f1; // ω147: 1.38336003

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd296; ram_i_data1 = 32'h401a964f; // θ148: 2.41542411
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd297; ram_i_data1 = 32'hbff8962a; // ω148:-1.94208264

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd298; ram_i_data1 = 32'h401d6306; // θ149: 2.45916891
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd299; ram_i_data1 = 32'h40122b01; // ω149: 2.28387475

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd300; ram_i_data1 = 32'h3e6f7b20; // θ150: 0.23386812
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd301; ram_i_data1 = 32'hbfed90cb; // ω150:-1.85598123

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd302; ram_i_data1 = 32'hbfaf1bf3; // θ151:-1.36804044
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd303; ram_i_data1 = 32'h40114f55; // ω151: 2.27046704

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd304; ram_i_data1 = 32'h4009f94a; // θ152: 2.15584040
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd305; ram_i_data1 = 32'hbff649e7; // ω152:-1.92413032

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd306; ram_i_data1 = 32'hbfe85004; // θ153:-1.81494188
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd307; ram_i_data1 = 32'hbfeada08; // ω153:-1.83477879

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd308; ram_i_data1 = 32'h3ffabf99; // θ154: 1.95897210
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd309; ram_i_data1 = 32'h3fa70798; // ω154: 1.30491924

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd310; ram_i_data1 = 32'hbf48f756; // θ155:-0.78502405
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd311; ram_i_data1 = 32'h3fd53903; // ω155: 1.66580236

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd312; ram_i_data1 = 32'hbfef28fc; // θ156:-1.86843824
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd313; ram_i_data1 = 32'h3faf1b4c; // ω156: 1.36802053

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd314; ram_i_data1 = 32'hc007297a; // θ157:-2.11190653
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd315; ram_i_data1 = 32'hc03e3ee3; // ω157:-2.97258830

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd316; ram_i_data1 = 32'h4012d2f1; // θ158: 2.29412484
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd317; ram_i_data1 = 32'hbe9a9c4f; // ω158:-0.30197379

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd318; ram_i_data1 = 32'hbf9ba645; // θ159:-1.21601164
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd319; ram_i_data1 = 32'hc0461be5; // ω159:-3.09545255

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd320; ram_i_data1 = 32'h3fb1214e; // θ160: 1.38382888
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd321; ram_i_data1 = 32'h402cbe09; // ω160: 2.69909883

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd322; ram_i_data1 = 32'h3fee8612; // θ161: 1.86346650
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd323; ram_i_data1 = 32'hbf0f1e06; // ω161:-0.55905187

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd324; ram_i_data1 = 32'h40024fbb; // θ162: 2.03611636
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd325; ram_i_data1 = 32'h3e45cf91; // ω162: 0.19317462

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd326; ram_i_data1 = 32'hbeb98f63; // θ163:-0.36242208
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd327; ram_i_data1 = 32'hc02e0676; // ω163:-2.71914434

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd328; ram_i_data1 = 32'hc03c50be; // θ164:-2.94242811
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd329; ram_i_data1 = 32'h3f168d40; // ω164: 0.58809280

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd330; ram_i_data1 = 32'hbda56b9d; // θ165:-0.08077166
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd331; ram_i_data1 = 32'h3f1939e4; // ω165: 0.59853959

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd332; ram_i_data1 = 32'h4047798b; // θ166: 3.11679339
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd333; ram_i_data1 = 32'hc04887f7; // ω166:-3.13329864

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd334; ram_i_data1 = 32'hc0405a67; // θ167:-3.00551772
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd335; ram_i_data1 = 32'h3fc69b9c; // ω167: 1.55162382

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd336; ram_i_data1 = 32'h3ffef4a1; // θ168: 1.99184048
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd337; ram_i_data1 = 32'hbfc884b2; // ω168:-1.56654954

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd338; ram_i_data1 = 32'hbff01805; // θ169:-1.87573302
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd339; ram_i_data1 = 32'h3fa08ec8; // ω169: 1.25435734

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd340; ram_i_data1 = 32'hc01bd391; // θ170:-2.43478799
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd341; ram_i_data1 = 32'h3fb420f3; // ω170: 1.40725553

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd342; ram_i_data1 = 32'h3f5534b8; // θ171: 0.83283567
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd343; ram_i_data1 = 32'hc01d1f93; // ω171:-2.45505214

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd344; ram_i_data1 = 32'h40082905; // θ172: 2.12750363
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd345; ram_i_data1 = 32'hc01ebdb5; // ω172:-2.48032880

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd346; ram_i_data1 = 32'h3fdeab1b; // θ173: 1.73959672
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd347; ram_i_data1 = 32'h3fb4ca41; // ω173: 1.41242230

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd348; ram_i_data1 = 32'hc03c7c0c; // θ174:-2.94507122
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd349; ram_i_data1 = 32'h3fcfb967; // ω174: 1.62284553

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd350; ram_i_data1 = 32'hc00a1dc6; // θ175:-2.15806723
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd351; ram_i_data1 = 32'h3f93aa74; // ω175: 1.15363932

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd352; ram_i_data1 = 32'h3fc6295c; // θ176: 1.54813719
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd353; ram_i_data1 = 32'hbfe86d4b; // ω176:-1.81583536

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd354; ram_i_data1 = 32'h3f0f1170; // θ177: 0.55885983
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd355; ram_i_data1 = 32'h4041b0e7; // ω177: 3.02642226

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd356; ram_i_data1 = 32'h4044b8cb; // θ178: 3.07377887
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd357; ram_i_data1 = 32'h3f0c7670; // ω178: 0.54868221

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd358; ram_i_data1 = 32'h40328326; // θ179: 2.78925467
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd359; ram_i_data1 = 32'h3f46af9e; // ω179: 0.77611721

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd360; ram_i_data1 = 32'hbe75b510; // θ180:-0.23994851
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd361; ram_i_data1 = 32'h3ec38906; // ω180: 0.38190478

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd362; ram_i_data1 = 32'hc01c71a5; // θ181:-2.44443631
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd363; ram_i_data1 = 32'hbeba150c; // ω181:-0.36344182

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd364; ram_i_data1 = 32'hbe9d11d0; // θ182:-0.30677652
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd365; ram_i_data1 = 32'h40222b11; // ω182: 2.53387856

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd366; ram_i_data1 = 32'hbe6f1087; // θ183:-0.23346148
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd367; ram_i_data1 = 32'h3f6c2138; // ω183: 0.92238188

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd368; ram_i_data1 = 32'hc01a3e8a; // θ184:-2.41006708
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd369; ram_i_data1 = 32'hbfd87aef; // ω184:-1.69125164

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd370; ram_i_data1 = 32'h4027105b; // θ185: 2.61037326
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd371; ram_i_data1 = 32'h3df486d9; // ω185: 0.11939783

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd372; ram_i_data1 = 32'hc011180d; // θ186:-2.26709294
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd373; ram_i_data1 = 32'h400c89f6; // ω186: 2.19592047

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd374; ram_i_data1 = 32'hbfed2a5a; // θ187:-1.85285497
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd375; ram_i_data1 = 32'h3ec65de4; // ω187: 0.38743508

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd376; ram_i_data1 = 32'hc032a3cc; // θ188:-2.79124737
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd377; ram_i_data1 = 32'h3e8b4ead; // ω188: 0.27208462

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd378; ram_i_data1 = 32'h3e31d1b8; // θ189: 0.17365158
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd379; ram_i_data1 = 32'h3fb74aef; // ω189: 1.43197429

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd380; ram_i_data1 = 32'h4003184a; // θ190: 2.04835749
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd381; ram_i_data1 = 32'h3f8471a1; // ω190: 1.03471768

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd382; ram_i_data1 = 32'hbde6e5b3; // θ191:-0.11274280
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd383; ram_i_data1 = 32'hbf414610; // ω191:-0.75497532

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h3f2720aa; // action0:  0.65284216
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3fca6536; // action1:  1.58121371
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'hbffa6791; // action2: -1.95628560
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'hbf2d47c2; // action3: -0.67687619
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3ec5437d; // action4:  0.38528052
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbfd6a184; // action5: -1.67680407
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3fcb371e; // action6:  1.58761954
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbfecd69c; // action7: -1.85029936
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h3ff257b8; // action8:  1.89330196
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbfa242e4; // action9: -1.26766634
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h3ff49890; // action10:  1.91090584
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbf8cdd93; // action11: -1.10051191
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h3f50c4ef; // action12:  0.81550497
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h3f4995de; // action13:  0.78744304
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h3fc3218f; // action14:  1.52446163
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'hbe71b0c6; // action15: -0.23602590
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h3e6d1001; // action16:  0.23150636
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'hbf7c8489; // action17: -0.98639733
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'hbfb5a07a; // action18: -1.41895986
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h3fd6d937; // action19:  1.67850387
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'hbd636774; // action20: -0.05551858
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h3fa660d9; // action21:  1.29983056
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'hbf9dce57; // action22: -1.23285949
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbf54945f; // action23: -0.83038896
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbfaf9193; // action24: -1.37163007
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'hbffe9dd6; // action25: -1.98919177
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h3e9753ce; // action26:  0.29556125
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3eac4aa3; // action27:  0.33650693
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3e8edac7; // action28:  0.27901289
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbe9565bf; // action29: -0.29179189
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3ffc6c14; // action30:  1.97204828
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h3fc38018; // action31:  1.52734661
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h3fdc0f4d; // action32:  1.71921694
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'hbfe8935b; // action33: -1.81699693
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'hbecf9960; // action34: -0.40546703
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3f277b7d; // action35:  0.65422803
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'hbfb8b3f8; // action36: -1.44299221
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h3e00060e; // action37:  0.12502310
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbfa20975; // action38: -1.26591361
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h3f7107a7; // action39:  0.94152302
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'hbecfcc06; // action40: -0.40585345
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h3e1dc9c9; // action41:  0.15409006
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'hbf9fd892; // action42: -1.24879670
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbea5f61f; // action43: -0.32414338
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'hbfbdd41c; // action44: -1.48303556
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3fa68afb; // action45:  1.30111635
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbf39cd41; // action46: -0.72578818
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3fd70caa; // action47:  1.68007398
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h3ffd7866; // action48:  1.98023677
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h3f9ac734; // action49:  1.20920420
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbfb8f394; // action50: -1.44493341
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbfffd4d1; // action51: -1.99868214
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h3eaa8a9b; // action52:  0.33308873
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'hbed700f6; // action53: -0.41992921
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'hbf54e12d; // action54: -0.83156091
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'hbf97d84f; // action55: -1.18628871
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'hbfda7366; // action56: -1.70664668
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbf685604; // action57: -0.90756249
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3fe86d34; // action58:  1.81583261
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'hbda2b3d3; // action59: -0.07944455
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbf440eb7; // action60: -0.76584953
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3f8d997b; // action61:  1.10624635
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3dfbec74; // action62:  0.12300959
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3fa5c69b; // action63:  1.29512346
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'hbfa072a6; // action64: -1.25349879
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3fe762ba; // action65:  1.80770040
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h3ea5b235; // action66:  0.32362524
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbffa302a; // action67: -1.95459485
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3a9b932f; // action68:  0.00118694
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'hbfe20275; // action69: -1.76569998
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h3f450ea0; // action70:  0.76975441
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3ee2798d; // action71:  0.44233361
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'hbecc12fc; // action72: -0.39858234
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'hbe5d0b9c; // action73: -0.21586460
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'hbe82b6f6; // action74: -0.25530213
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'hbf758a3d; // action75: -0.95914060
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'hbf880b51; // action76: -1.06284535
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h3e92c59a; // action77:  0.28666383
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbfd35f98; // action78: -1.65135479
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbf43c524; // action79: -0.76472688
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3fc66595; // action80:  1.54997504
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3ee608c1; // action81:  0.44928554
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'hbf3dbcd9; // action82: -0.74116284
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'hbf8e0a79; // action83: -1.10969460
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbf380216; // action84: -0.71878183
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbf9d7a9d; // action85: -1.23030436
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h3f7d6881; // action86:  0.98987585
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3f8f01a9; // action87:  1.11723816
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h3fc019da; // action88:  1.50078893
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbfa2c782; // action89: -1.27171350
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3fcc5241; // action90:  1.59626019
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3fc2e832; // action91:  1.52271104
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbf83fbf7; // action92: -1.03112686
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'hbfec01f7; // action93: -1.84380996
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3f9a3ad2; // action94:  1.20492005
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h3f1c3f11; // action95:  0.61033732
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'hbf749a8c; // action96: -0.95548320
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3f93a925; // action97:  1.15359938
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbf161003; // action98: -0.58618182
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3f1b8f95; // action99:  0.60765964
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h3d8a75ce; // action100:  0.06760751
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'hbf019bb9; // action101: -0.50628239
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3feb8977; // action102:  1.84013259
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbf1d68b2; // action103: -0.61487877
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h3fe786a9; // action104:  1.80879700
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbf5261af; // action105: -0.82180303
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3f030200; // action106:  0.51174927
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbfa018cc; // action107: -1.25075674
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3f8ac944; // action108:  1.08426714
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'hbf19a0da; // action109: -0.60011065
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'hbf6d2404; // action110: -0.92633080
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbfb28cc7; // action111: -1.39492118
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3d03c691; // action112:  0.03217179
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h3f6597d5; // action113:  0.89684802
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h3fe69819; // action114:  1.80151665
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3fd53005; // action115:  1.66552794
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3fa8dfec; // action116:  1.31933355
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'hbec8ddd9; // action117: -0.39231756
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'hbf6e4f29; // action118: -0.93089539
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'hbf350229; // action119: -0.70706421
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'hbf393c3c; // action120: -0.72357535
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3f183071; // action121:  0.59448916
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h3fd92961; // action122:  1.69657528
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3fecbdfc; // action123:  1.84954786
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3f6ee802; // action124:  0.93322766
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h3db91f1d; // action125:  0.09039138
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbfe0da0b; // action126: -1.75665414
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3f98e079; // action127:  1.19435036
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'hbf03a9da; // action128: -0.51431048
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3fec6031; // action129:  1.84668553
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'hbfbf90f0; // action130: -1.49661064
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h3f60e5f0; // action131:  0.87850857
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'hbf50004b; // action132: -0.81250447
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3f2c3cd9; // action133:  0.67280346
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3fb040f3; // action134:  1.37698209
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h3f76650d; // action135:  0.96247941
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h3e63c523; // action136:  0.22243170
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'hbf8b228d; // action137: -1.08699191
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h3fc20965; // action138:  1.51591170
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h3ee79f10; // action139:  0.45238543
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'hbfc7c607; // action140: -1.56073081
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'hbd733fba; // action141: -0.05938695
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'hbf4287d6; // action142: -0.75988519
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h3fa38398; // action143:  1.27745342
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3ede07f5; // action144:  0.43365446
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h3ed56bf2; // action145:  0.41683918
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'hbea80e01; // action146: -0.32823184
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h3e941098; // action147:  0.28918910
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3f82d9f4; // action148:  1.02227640
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbf8c74c7; // action149: -1.09731376
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'hbf1ba77c; // action150: -0.60802436
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbfdfeb17; // action151: -1.74936187
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3f8535b5; // action152:  1.04070151
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3fd7cbd0; // action153:  1.68590736
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'hbfcb88c4; // action154: -1.59011126
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h3f4720bd; // action155:  0.77784330
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbea5c336; // action156: -0.32375497
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h3fc93aab; // action157:  1.57210290
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbf72220f; // action158: -0.94583219
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h3f60415c; // action159:  0.87599730
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbfcaa70f; // action160: -1.58322322
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'hbfc7f274; // action161: -1.56208658
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h3fc775a9; // action162:  1.55827820
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h3fa09651; // action163:  1.25458729
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h3f8e951a; // action164:  1.11392522
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'hbeebfc60; // action165: -0.46090984
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbfb7a093; // action166: -1.43458784
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbfa217c8; // action167: -1.26635075
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3fba6dae; // action168:  1.45647216
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h3f080fbc; // action169:  0.53149009
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbfb23fb6; // action170: -1.39256930
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3fb6363f; // action171:  1.42353046
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3f0b99aa; // action172:  0.54531348
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3ec82b5a; // action173:  0.39095575
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3d98fd62; // action174:  0.07470204
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'hbf914adf; // action175: -1.13509738
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3ffc71b3; // action176:  1.97221982
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h3fd1ad78; // action177:  1.63810635
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h3e6c7fde; // action178:  0.23095652
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbee0643d; // action179: -0.43826476
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'hbff8131e; // action180: -1.93808341
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h3fd5e872; // action181:  1.67115617
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbfcbd336; // action182: -1.59238315
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h3e53fe8a; // action183:  0.20702568
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3f99d45f; // action184:  1.20179355
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h3fa2a212; // action185:  1.27057099
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3fb211b0; // action186:  1.39116478
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'hbff93797; // action187: -1.94700897
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbf7a8d1c; // action188: -0.97871566
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbf797547; // action189: -0.97444576
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h3d09cd3f; // action190:  0.03364300
            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h3e65938f; // action191:  0.22419570

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd2; new_round = 1'b1; // clear flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 1:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbffef6aa; // action0: -1.99190259
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3ea41cb4; // action1:  0.32053149
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'hbfaa5e93; // action2: -1.33101118
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3f12fcd3; // action3:  0.57417029
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'hbea1dcde; // action4: -0.31613821
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h3fae63ab; // action5:  1.36241663
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'hbfd682ef; // action6: -1.67587078
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbfd796c6; // action7: -1.68428874
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h3ff8fe5e; // action8:  1.94526267
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h3fe889c2; // action9:  1.81670403
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h3fef31ab; // action10:  1.86870325
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbfa7e621; // action11: -1.31171048
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'hbf2cb47b; // action12: -0.67462891
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h3ec8e9d6; // action13:  0.39240903
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h3ee6b103; // action14:  0.45056924
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3fb18b5c; // action15:  1.38706541
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h3feaf3c1; // action16:  1.83556378
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h3fc34409; // action17:  1.52551377
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h3f6a3e65; // action18:  0.91501456
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h3f8596ea; // action19:  1.04366803
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h3e27abb4; // action20:  0.16374093
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h3ec95a71; // action21:  0.39326814
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h3f066f70; // action22:  0.52513790
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbfe0b1d0; // action23: -1.75542641
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbe0c4d87; // action24: -0.13701449
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3f89b9ce; // action25:  1.07598281
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'hbf821162; // action26: -1.01615548
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3fa5c090; // action27:  1.29493904
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3ffde62a; // action28:  1.98358655
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h3e0b6d6a; // action29:  0.13615957
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3f877221; // action30:  1.05817044
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbfdfd60a; // action31: -1.74871945
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h3e4b8632; // action32:  0.19875410
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'hbe80c4e1; // action33: -0.25150207
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'hbfcfb8f0; // action34: -1.62283134
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3fb41615; // action35:  1.40692389
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3f30d5b8; // action36:  0.69076109
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'hbff7f1ec; // action37: -1.93707037
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbfcd6eda; // action38: -1.60494542
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'hbfb976a7; // action39: -1.44893348
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3ffd4558; // action40:  1.97867870
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h3e80c91b; // action41:  0.25153431
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3ff660e8; // action42:  1.92483234
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h3e0b0389; // action43:  0.13575567
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3e713e99; // action44:  0.23559035
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3f0d410d; // action45:  0.55177385
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbfe8d4f6; // action46: -1.81899905
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3dbfb040; // action47:  0.09359789
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h3fb753cd; // action48:  1.43224490
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h3e389dbf; // action49:  0.18028925
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbfa28919; // action50: -1.26980889
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbf1a6264; // action51: -0.60306382
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbfb24f36; // action52: -1.39304233
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'hbe9fb0cc; // action53: -0.31189573
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3f5e5494; // action54:  0.86847806
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h3f7827bd; // action55:  0.96935636
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h3fefa3d6; // action56:  1.87218738
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h3dc9bd90; // action57:  0.09850609
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'hbf82c257; // action58: -1.02155578
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h3fc2eafc; // action59:  1.52279615
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbfe450bf; // action60: -1.78371418
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'hbeb4d1c6; // action61: -0.35316294
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3e315970; // action62:  0.17319274
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'hbfccd2af; // action63: -1.60017955
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3ff23bc5; // action64:  1.89244902
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3f7fe7cd; // action65:  0.99963075
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h3f25b52d; // action66:  0.64729577
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h3da43f78; // action67:  0.08019918
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3fdd016e; // action68:  1.72660613
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3f824b1c; // action69:  1.01791716
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h3f6ad9a2; // action70:  0.91738331
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'hbf6237c0; // action71: -0.88366318
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3baee419; // action72:  0.00533725
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'hbef85b78; // action73: -0.48507285
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'hbe9ce261; // action74: -0.30641463
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3fd64799; // action75:  1.67405999
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'hbfa4362c; // action76: -1.28290319
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbe693c40; // action77: -0.22776890
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbf62d568; // action78: -0.88606882
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbff97120; // action79: -1.94876480
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3e6957dd; // action80:  0.22787423
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'hbf053ce4; // action81: -0.52046037
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'hbfa8d0bf; // action82: -1.31887043
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'hbf311c53; // action83: -0.69183844
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h3f35542d; // action84:  0.70831567
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbfa81941; // action85: -1.31327069
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h3faa6782; // action86:  1.33128381
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'hbf2f485a; // action87: -0.68469775
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h3f887e0f; // action88:  1.06634700
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbe5499f7; // action89: -0.20761858
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3f6a5fce; // action90:  0.91552436
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3b244d27; // action91:  0.00250704
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h3fb79b88; // action92:  1.43443394
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'hbf313822; // action93: -0.69226277
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3f547b89; // action94:  0.83001000
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'hbf920f3f; // action95: -1.14109027
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h3dca562d; // action96:  0.09879718
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'hbfc6c2e9; // action97: -1.55282319
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbf4cfeb6; // action98: -0.80076158
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3fe9990d; // action99:  1.82498324
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'hbf7120ef; // action100: -0.94190878
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'hbfe30417; // action101: -1.77356231
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'hbff6128c; // action102: -1.92244101
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h3fc4f694; // action103:  1.53877497
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'hbf880a4a; // action104: -1.06281400
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbf33c3b8; // action105: -0.70220518
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3f96f486; // action106:  1.17933726
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h3ff896d7; // action107:  1.94210327
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3e0414b5; // action108:  0.12898524
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'hbe853a8c; // action109: -0.26021230
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'hbfdfb4e2; // action110: -1.74770761
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h3f24c8ee; // action111:  0.64369094
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'hbfb7856b; // action112: -1.43375909
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'hbeee6da1; // action113: -0.46568015
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'hbf99bb52; // action114: -1.20102906
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3ef18437; // action115:  0.47171184
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3fc4c25b; // action116:  1.53718126
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3fe7a604; // action117:  1.80975389
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3ff62564; // action118:  1.92301607
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'hbfa32144; // action119: -1.27445269
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'hbfe318a7; // action120: -1.77418983
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3f99a9a0; // action121:  1.20048904
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h3fc82310; // action122:  1.56357002
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3f83ba0f; // action123:  1.02911556
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3fd2f98b; // action124:  1.64824045
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h3fd29657; // action125:  1.64521301
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h3f734ca7; // action126:  0.95038837
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'hbfefd414; // action127: -1.87365961
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h3fbbeb13; // action128:  1.46811140
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3fbffd3e; // action129:  1.49991584
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h3ff242e5; // action130:  1.89266646
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbfc45ebc; // action131: -1.53414106
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'hbf9953c9; // action132: -1.19786942
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'hbf573e76; // action133: -0.84079683
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'hbf65261b; // action134: -0.89511269
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'hbf98c3a2; // action135: -1.19347024
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'hbfe7f24d; // action136: -1.81208193
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'hbff4af2e; // action137: -1.91159606
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h3fff57ae; // action138:  1.99486327
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'hbffcb0b6; // action139: -1.97414279
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'hbfc12d9b; // action140: -1.50920427
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'hbfb52385; // action141: -1.41514647
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'hbfec7885; // action142: -1.84742796
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'hbfee2c8a; // action143: -1.86073422
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3fedf7f8; // action144:  1.85912991
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h3f691053; // action145:  0.91040534
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h3fab87cd; // action146:  1.34008181
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbf102da1; // action147: -0.56319624
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3ff52f6f; // action148:  1.91551006
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbfbd4f5c; // action149: -1.47898436
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'hbfe73c25; // action150: -1.80652297
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbf7dff3a; // action151: -0.99217570
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'hbf34d529; // action152: -0.70637757
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3f3a0a24; // action153:  0.72671723
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h3e7cf899; // action154:  0.24704207
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h3f75f7c3; // action155:  0.96081179
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h3cbf015d; // action156:  0.02331608
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbf0ca6b0; // action157: -0.54941845
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbf2e5713; // action158: -0.68101615
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h3ffd9091; // action159:  1.98097432
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbff6666f; // action160: -1.92500103
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'hbf82266a; // action161: -1.01679730
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h3fdd1126; // action162:  1.72708583
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h3f4f4701; // action163:  0.80967718
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbed1a4fd; // action164: -0.40946189
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'hbfd4d134; // action165: -1.66263437
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h3f16ce89; // action166:  0.58908898
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbf0cb7b7; // action167: -0.54967827
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3fd90571; // action168:  1.69547856
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbe74b958; // action169: -0.23898828
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbfaec6a4; // action170: -1.36543703
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3e32e577; // action171:  0.17470346
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'hbff3eed7; // action172: -1.90572631
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3eb9535c; // action173:  0.36196411
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3fc80ab6; // action174:  1.56282687
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'hbf860174; // action175: -1.04691935
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3f2409d7; // action176:  0.64077514
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'hbf5444e7; // action177: -0.82917637
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbf1256eb; // action178: -0.57163876
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbff88f64; // action179: -1.94187593
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'hbf940a32; // action180: -1.15656114
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h3f6e0793; // action181:  0.92980307
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbfa12da2; // action182: -1.25920510
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'hbfa52b5f; // action183: -1.29038608
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'hbec608c7; // action184: -0.38678572
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h3f97f033; // action185:  1.18701780
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3e154946; // action186:  0.14578733
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'hbf709198; // action187: -0.93972158
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbfdbaa6d; // action188: -1.71613848
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbdd35097; // action189: -0.10318106
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'hbdd21c97; // action190: -0.10259359
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'hbffc5c30; // action191: -1.97156334

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 2:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbe6761a1; // action0: -0.22595836
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3ff225f1; // action1:  1.89178288
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3fa1c6fd; // action2:  1.26388514
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3e929b78; // action3:  0.28634238
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3f376f20; // action4:  0.71653938
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbfaa3eb3; // action5: -1.33003843
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3ec2012e; // action6:  0.37891525
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbfab16cf; // action7: -1.33663356
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'hbf096046; // action8: -0.53662527
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbffd5fdc; // action9: -1.97948790
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'hbf0a94e7; // action10: -0.54133457
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h3db86bd5; // action11:  0.09004942
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h3fcabeef; // action12:  1.58395183
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbfb1d267; // action13: -1.38923347
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbfb764fc; // action14: -1.43276930
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3f2d7901; // action15:  0.67762762
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'hbf2ed8fe; // action16: -0.68299854
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'hbeb0d8ee; // action17: -0.34540504
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h3f7058c1; // action18:  0.93885428
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbfc1e241; // action19: -1.51471722
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h3ea413c0; // action20:  0.32046318
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbe80b2a6; // action21: -0.25136298
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h3fc16153; // action22:  1.51078260
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h3f66b078; // action23:  0.90113020
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbee77dbf; // action24: -0.45213124
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3fba335d; // action25:  1.45469248
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'hbeea8e19; // action26: -0.45811537
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3fc03929; // action27:  1.50174439
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'hbee85e4a; // action28: -0.45384437
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h3f147438; // action29:  0.57989836
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3f8ded3a; // action30:  1.10880208
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h3fe1d826; // action31:  1.76440883
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbfe4e1df; // action32: -1.78814304
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'hbee28652; // action33: -0.44243103
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'hbf1f9086; // action34: -0.62329900
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3ca560f8; // action35:  0.02018784
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3eea7359; // action36:  0.45791128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'hbfec6f29; // action37: -1.84714234
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h3f57ce8e; // action38:  0.84299552
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'hbfcae3b8; // action39: -1.58507442
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3f2ca2c3; // action40:  0.67435855
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h3f3ae2a3; // action41:  0.73002070
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3f4f5bdc; // action42:  0.80999541
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbfd7e43a; // action43: -1.68665242
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'hbf03b443; // action44: -0.51446933
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'hbf259e0c; // action45: -0.64694285
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbfaadaae; // action46: -1.33479857
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3f38a58a; // action47:  0.72127593
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h3fb183ab; // action48:  1.38683069
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbfefcebf; // action49: -1.87349689
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbfe46506; // action50: -1.78433299
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbfe56dac; // action51: -1.79240942
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbf714149; // action52: -0.94240242
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h3f993ffa; // action53:  1.19726491
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3e479ae7; // action54:  0.19492684
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'hbfaf7e20; // action55: -1.37103653
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h3f07ff9c; // action56:  0.53124404
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h3f1d5c46; // action57:  0.61468923
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'hbe8c7232; // action58: -0.27430874
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'hbff4f2b6; // action59: -1.91365695
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbe93ce21; // action60: -0.28868201
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3ebb16a3; // action61:  0.36540708
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'hbd9c5f6e; // action62: -0.07635389
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3ee6efac; // action63:  0.45104730
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'hbf95c77c; // action64: -1.17015028
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3fd18b9a; // action65:  1.63707280
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h3fe4c207; // action66:  1.78717124
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbff6afe5; // action67: -1.92724288
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'hbff8ed4f; // action68: -1.94474208
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'hbfa30577; // action69: -1.27360427
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'hbfe77e80; // action70: -1.80854797
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'hbf81e389; // action71: -1.01475632
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'hbf9a7c74; // action72: -1.20692301
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3fa8060c; // action73:  1.31268454
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3e8a661a; // action74:  0.27031022
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'hbf097922; // action75: -0.53700459
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h3eb38386; // action76:  0.35061282
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h3f166b12; // action77:  0.58757126
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbec6573c; // action78: -0.38738430
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbf13ef4d; // action79: -0.57787019
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'hbf1da69a; // action80: -0.61582339
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3f46064c; // action81:  0.77353358
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h3dc4e791; // action82:  0.09614480
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h3fb53cd2; // action83:  1.41591859
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbf935511; // action84: -1.15103352
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h3ff8c6c5; // action85:  1.94356596
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'hbf9871f4; // action86: -1.19097757
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3feff664; // action87:  1.87470675
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbfff174d; // action88: -1.99289858
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbe10fd22; // action89: -0.14159063
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'hbfcb6982; // action90: -1.58915734
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3e03826d; // action91:  0.12842722
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbf8fdc1d; // action92: -1.12390482
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h3eb0cb48; // action93:  0.34530091
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3ef5ff26; // action94:  0.48046225
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'hbf89c2d4; // action95: -1.07625818
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'hbe3d7b9f; // action96: -0.18504189
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3f131bf2; // action97:  0.57464516
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbf6e6cbc; // action98: -0.93134665
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3faff4e2; // action99:  1.37466073
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h3f8a4413; // action100:  1.08020246
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h3d91a083; // action101:  0.07110693
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3fd9cc3d; // action102:  1.70154536
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h3f34dd06; // action103:  0.70649755
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'hbe1e5bdb; // action104: -0.15464728
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h3fae0bba; // action105:  1.35973287
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3f685da8; // action106:  0.90767908
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbf59b859; // action107: -0.85046917
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3eaa9e9b; // action108:  0.33324131
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3ec656ee; // action109:  0.38738197
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'hbf9f019d; // action110: -1.24223673
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbfe12e92; // action111: -1.75923371
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3c0153c8; // action112:  0.00789351
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h3f88dc18; // action113:  1.06921673
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h3fbb7797; // action114:  1.46458709
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'hbfc2c602; // action115: -1.52166772
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3eea7024; // action116:  0.45788682
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'hbe8b9fad; // action117: -0.27270260
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3fe1a0ca; // action118:  1.76271939
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3fb3ce96; // action119:  1.40474200
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'hbf340c09; // action120: -0.70330864
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3f872455; // action121:  1.05579627
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h3faeb301; // action122:  1.36483777
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'hbf28b445; // action123: -0.65900069
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3eccfb4f; // action124:  0.40035483
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h3fe1444e; // action125:  1.75989699
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbf464ed7; // action126: -0.77464050
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3fc8889f; // action127:  1.56666934
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'hbf4f6dba; // action128: -0.81026804
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'hbec7b42e; // action129: -0.39004654
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h3fcf1b07; // action130:  1.61801231
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbf6771e7; // action131: -0.90408176
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'hbfd10f7c; // action132: -1.63328505
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'hbff1bb00; // action133: -1.88851929
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'hbfa18a96; // action134: -1.26204181
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h3f4dc1b4; // action135:  0.80373693
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'hbfb014ae; // action136: -1.37563109
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'hbfb2e450; // action137: -1.39759254
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h3fd51b7a; // action138:  1.66490102
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h3f9671f9; // action139:  1.17535317
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h3fabe8a2; // action140:  1.34303689
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'hbf6ceeb0; // action141: -0.92551708
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'hbf0eeced; // action142: -0.55830270
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'hbf2acd85; // action143: -0.66719848
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3e89cf4b; // action144:  0.26915964
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'hbfcb3bf0; // action145: -1.58776665
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'hbf33ae3e; // action146: -0.70187747
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbf295b65; // action147: -0.66155082
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3ed2c0f0; // action148:  0.41162825
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbe125a36; // action149: -0.14292225
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'hbebb2176; // action150: -0.36548966
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h3f35b0b0; // action151:  0.70972729
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'hbff9027d; // action152: -1.94538844
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3f9961be; // action153:  1.19829535
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'hbeccfc31; // action154: -0.40036157
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h3f67bceb; // action155:  0.90522641
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbfe8bc9c; // action156: -1.81825590
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbf804974; // action157: -1.00224161
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h3f746278; // action158:  0.95462751
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'hbffbbaa1; // action159: -1.96663296
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbfda6184; // action160: -1.70610094
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h3f86c527; // action161:  1.05289161
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h3f962cb8; // action162:  1.17323971
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h3fc10dfd; // action163:  1.50823939
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbf88d156; // action164: -1.06888843
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'hbf951c40; // action165: -1.16492462
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbfd2282b; // action166: -1.64185083
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h3e604af0; // action167:  0.21903586
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3ff82c5c; // action168:  1.93885374
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbfcbc3e8; // action169: -1.59191608
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h3dcdd8d6; // action170:  0.10051124
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3fab1194; // action171:  1.33647394
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'hbf3d7c63; // action172: -0.74017924
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'hbfe344d4; // action173: -1.77553797
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3e3cefd6; // action174:  0.18450865
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3f9132e8; // action175:  1.13436604
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'hbfc39ca3; // action176: -1.52821767
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h3fc385ba; // action177:  1.52751851
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h3ee0d977; // action178:  0.43915913
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h3f8034a6; // action179:  1.00160670
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'hbf53c228; // action180: -0.82718134
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbfd11e5a; // action181: -1.63373876
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbe1cb322; // action182: -0.15302709
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h3e316d0a; // action183:  0.17326751
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'hbf8730bf; // action184: -1.05617511
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbd506d99; // action185: -0.05088577
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3fa93be0; // action186:  1.32213974
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'hbfbd9080; // action187: -1.48097229
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbf966d9f; // action188: -1.17522037
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h3c14e225; // action189:  0.00908712
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'hbf0878c6; // action190: -0.53309286
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'hbef60051; // action191: -0.48047116

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 3:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbf8f23c6; // action0: -1.11827922
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'hbfbc16f2; // action1: -1.46945024
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3e0860af; // action2:  0.13318132
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3f37ea2a; // action3:  0.71841681
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3fb4f572; // action4:  1.41374040
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbf0ab314; // action5: -0.54179502
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'hbd4fc47e; // action6: -0.05072450
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h3e14bb64; // action7:  0.14524609
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'hbf1e8429; // action8: -0.61920410
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbf8aa3df; // action9: -1.08312595
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'hbf6aaf94; // action10: -0.91674161
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbfc96111; // action11: -1.57327473
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h3f100441; // action12:  0.56256491
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbfa5fbfc; // action13: -1.29675245
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbf0a4a9b; // action14: -0.54020089
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3faaa82e; // action15:  1.33325744
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'hbf6f8fb0; // action16: -0.93578625
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h3fd9a856; // action17:  1.70044971
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h3fbd6cf5; // action18:  1.47988760
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbf5a1986; // action19: -0.85195196
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h3fbd10d6; // action20:  1.47707629
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbfda66d3; // action21: -1.70626295
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'hbfca6597; // action22: -1.58122528
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h3fe5aa72; // action23:  1.79426408
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h3ebaf299; // action24:  0.36513212
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'hbfc3937d; // action25: -1.52793849
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h3d8f1c6d; // action26:  0.06987844
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3e0ee14a; // action27:  0.13953128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3fb40345; // action28:  1.40634978
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h3eb93880; // action29:  0.36175919
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'hbf5d5733; // action30: -0.86461180
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbf8947d9; // action31: -1.07250512
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h3f13fec2; // action32:  0.57810605
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3f82e8b1; // action33:  1.02272618
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'hbe9de628; // action34: -0.30839658
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'hbd7cf27f; // action35: -0.06175470
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3f2a6bdc; // action36:  0.66570830
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h3fa7f442; // action37:  1.31214166
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbff52a2a; // action38: -1.91534925
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h3f89f1a6; // action39:  1.07768703
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'hbe6a1305; // action40: -0.22858818
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbee2ab93; // action41: -0.44271526
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'hbfc259db; // action42: -1.51836717
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbf6ff2e1; // action43: -0.93729979
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'hbf41dfe1; // action44: -0.75732237
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3f3686ae; // action45:  0.71299255
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbf26118c; // action46: -0.64870524
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3f9a6809; // action47:  1.20629990
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'hbfc05c5d; // action48: -1.50281870
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbfe4b769; // action49: -1.78684723
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbf74b666; // action50: -0.95590818
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h3f466143; // action51:  0.77492160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbfa03e58; // action52: -1.25190258
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'hbf886851; // action53: -1.06568348
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3de3d50b; // action54:  0.11124619
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h3fbbcd7b; // action55:  1.46720827
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'hbf783a41; // action56: -0.96963888
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h3f5decfc; // action57:  0.86689734
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3f124746; // action58:  0.57140005
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h3f8c9d87; // action59:  1.09855735
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbf494688; // action60: -0.78623247
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3fb3f20b; // action61:  1.40582407
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3e2fbd43; // action62:  0.17162041
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3fa038c2; // action63:  1.25173211
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3f476905; // action64:  0.77894622
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'hbda5aaa8; // action65: -0.08089191
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbffe3a35; // action66: -1.98615134
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h3ee9a7e5; // action67:  0.45635906
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3fd3e7ab; // action68:  1.65550745
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3f4257e8; // action69:  0.75915384
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'hbe2efaa1; // action70: -0.17087795
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3f7dd059; // action71:  0.99146038
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3e186f3d; // action72:  0.14886184
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3f9a4a52; // action73:  1.20539308
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3efbb134; // action74:  0.49158633
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3f83334c; // action75:  1.02500296
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'hbe4d0e50; // action76: -0.20024991
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbfc53745; // action77: -1.54074919
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h3e869c3e; // action78:  0.26291078
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbf8996ff; // action79: -1.07492054
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3ffc1100; // action80:  1.96926880
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3fc4eb8c; // action81:  1.53843832
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h3fa91080; // action82:  1.32081604
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'hbd562cc5; // action83: -0.05228879
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbff2ebb7; // action84: -1.89781845
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbf0348e1; // action85: -0.51283079
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'hbf8e6c34; // action86: -1.11267710
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3ffb4e76; // action87:  1.96333194
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbfd12e99; // action88: -1.63423455
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbf387c9b; // action89: -0.72065133
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3f48d043; // action90:  0.78442782
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3f4e29d8; // action91:  0.80532598
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h3f178d84; // action92:  0.59200311
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'hbef70e49; // action93: -0.48253086
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'hbf85f79f; // action94: -1.04661930
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h3f9a849d; // action95:  1.20717204
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h3fc0e7dc; // action96:  1.50707579
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3fa3b67a; // action97:  1.27900624
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbf8bd50f; // action98: -1.09243953
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'hbfe7e479; // action99: -1.81165993
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h3f4e08cb; // action100:  0.80482167
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'hbee17c73; // action101: -0.44040260
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'hbfdb62d9; // action102: -1.71395409
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbb91ec67; // action103: -0.00445323
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h3f8fe3c7; // action104:  1.12413871
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h3f3207c0; // action105:  0.69543076
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3f91f428; // action106:  1.14026356
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbf8d559a; // action107: -1.10417485
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3fb2628a; // action108:  1.39363217
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'hbf25f59c; // action109: -0.64827895
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h3fbbb12e; // action110:  1.46634459
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbfd87b1e; // action111: -1.69125724
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3f8d8ad0; // action112:  1.10579872
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'hbecb4177; // action113: -0.39698383
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'hbf9248f5; // action114: -1.14285147
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3eea3e94; // action115:  0.45750868
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3fcce105; // action116:  1.60061705
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'hbd8c6e54; // action117: -0.06856981
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3f35ad79; // action118:  0.70967823
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'hbf402b13; // action119: -0.75065726
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h3e172643; // action120:  0.14760689
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3fc1166b; // action121:  1.50849664
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h3fd5fca7; // action122:  1.67177284
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3f7c8194; // action123:  0.98635221
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3e022bd5; // action124:  0.12712033
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'hbf21029c; // action125: -0.62894607
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h3f091c5d; // action126:  0.53558904
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3fced0b7; // action127:  1.61574447
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h3f43d45d; // action128:  0.76495916
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'hbde70101; // action129: -0.11279488
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h3f58298e; // action130:  0.84438407
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbfa809b4; // action131: -1.31279612
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h3f673b29; // action132:  0.90324646
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3e37dc16; // action133:  0.17955050
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'hbcd03f2d; // action134: -0.02542075
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'hbf818e90; // action135: -1.01216316
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'hbf4211d3; // action136: -0.75808448
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'hbf1acc78; // action137: -0.60468245
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h3f5410ce; // action138:  0.82838142
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h3fd16e98; // action139:  1.63618755
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h3f97519f; // action140:  1.18217838
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h3f556f8e; // action141:  0.83373344
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3f7bc10e; // action142:  0.98341453
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'hbf4f241c; // action143: -0.80914474
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'hbf6746f2; // action144: -0.90342629
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h3ecdcaa9; // action145:  0.40193680
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h3faf3c87; // action146:  1.36903465
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h3f4f2fc1; // action147:  0.80932242
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3f3c4469; // action148:  0.73541886
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h3f9f8658; // action149:  1.24628735
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'hbfe3b9b9; // action150: -1.77910531
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbf1750b9; // action151: -0.59107548
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3d09982d; // action152:  0.03359239
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'hbddd4ca7; // action153: -0.10805636
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'hbff63922; // action154: -1.92361856
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h3edf20e9; // action155:  0.43579796
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h3fb513bd; // action156:  1.41466486
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbfe0e5cf; // action157: -1.75701320
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbfb65499; // action158: -1.42445672
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h3e42570c; // action159:  0.18978518
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h3f270eaf; // action160:  0.65256780
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'hbf924c1b; // action161: -1.14294755
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'hbda84c13; // action162: -0.08217635
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'hbfafbb14; // action163: -1.37289667
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbee4b3a2; // action164: -0.44668299
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3f956636; // action165:  1.16718173
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h3f244d1e; // action166:  0.64180171
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbe369940; // action167: -0.17831898
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'hbea7b35e; // action168: -0.32754034
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbe1c2c42; // action169: -0.15251258
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h3e61d6ee; // action170:  0.22054645
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'hbfa48d5f; // action171: -1.28556430
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'hbfb741ff; // action172: -1.43170154
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3f9d86c7; // action173:  1.23067558
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'hbf420743; // action174: -0.75792331
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3eaea648; // action175:  0.34111238
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'hbf0c65c9; // action176: -0.54842812
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'hbfd73777; // action177: -1.68138015
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbe8851fd; // action178: -0.26625052
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbfcc47e3; // action179: -1.59594381
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'hbde17c08; // action180: -0.11009985
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h3fa5959b; // action181:  1.29362810
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h3eb6eca8; // action182:  0.35727429
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h3f413e42; // action183:  0.75485623
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3e2c4d81; // action184:  0.16826440
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbf63faf9; // action185: -0.89054829
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3fe0871d; // action186:  1.75412333
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h3f86c3ca; // action187:  1.05285001
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbfaa7aff; // action188: -1.33187854
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbf3695dd; // action189: -0.71322423
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h3fbacb9c; // action190:  1.45933867
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h3e1cf1e4; // action191:  0.15326649

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 4:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbec2e077; // action0: -0.38061878
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3f1ef853; // action1:  0.62097663
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3fd64f21; // action2:  1.67428982
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'hbe403276; // action3: -0.18769249
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'hbf4cf9c2; // action4: -0.80068600
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbf561790; // action5: -0.83629704
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3f2da3da; // action6:  0.67828143
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbfa7278b; // action7: -1.30589426
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'hbefa3372; // action8: -0.48867375
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbfeb302c; // action9: -1.83740759
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h3fb08c51; // action10:  1.37928212
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbf236552; // action11: -0.63826478
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'hbf696542; // action12: -0.91170132
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbf0e2b87; // action13: -0.55535167
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h3f507bed; // action14:  0.81439096
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3f5b13b2; // action15:  0.85576928
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'hbea4d938; // action16: -0.32196975
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h3f6819ed; // action17:  0.90664560
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'hbeae0947; // action18: -0.33991453
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbfca8624; // action19: -1.58221865
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h3f3b6878; // action20:  0.73206282
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbf81b99e; // action21: -1.01347709
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'hbff3228f; // action22: -1.89949214
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbf5a753e; // action23: -0.85335147
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h3f1a012c; // action24:  0.60158038
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3da51449; // action25:  0.08060510
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'hbdab9842; // action26: -0.08378650
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3fac2180; // action27:  1.34477234
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3fddef51; // action28:  1.73386586
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h3fa4c3dd; // action29:  1.28722727
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3e558dbf; // action30:  0.20854853
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h3f0439d4; // action31:  0.51650739
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbed97f1f; // action32: -0.42479798
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'hbf853120; // action33: -1.04056168
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'hbf05c2bf; // action34: -0.52250284
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3f3bb959; // action35:  0.73329693
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'hbd7fda96; // action36: -0.06246432
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'hbf3dcd2d; // action37: -0.74141198
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbf3b8f8c; // action38: -0.73265910
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h3e046f81; // action39:  0.12933160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3ff0f2fc; // action40:  1.88241529
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbffcbb42; // action41: -1.97446465
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3fcfc60a; // action42:  1.62323117
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h3fba3a78; // action43:  1.45490932
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3f94d6ee; // action44:  1.16280913
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'hbd1a18a8; // action45: -0.03762117
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h3ec67c58; // action46:  0.38766742
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3e997d09; // action47:  0.29978207
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'hbf1f5e3e; // action48: -0.62253177
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbf72e96e; // action49: -0.94887435
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h3f933eb0; // action50:  1.15035057
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbf38659d; // action51: -0.72030050
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h3ea60812; // action52:  0.32428032
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'hbfa4df06; // action53: -1.28805614
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'hbf87c09e; // action54: -1.06056571
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h3f4d9bb3; // action55:  0.80315703
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'hbf924aab; // action56: -1.14290369
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbedeff67; // action57: -0.43554232
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'hbe090522; // action58: -0.13380864
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'hbf931e5c; // action59: -1.14936399
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbfac00f6; // action60: -1.34377933
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'hbe5c836c; // action61: -0.21534508
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3fdc17d6; // action62:  1.71947742
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'hbfac502e; // action63: -1.34619689
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'hbf20b238; // action64: -0.62771940
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3f8bd066; // action65:  1.09229732
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbfa84f40; // action66: -1.31491852
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h3f175f56; // action67:  0.59129846
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3fccefa1; // action68:  1.60106289
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3f1cadbc; // action69:  0.61202598
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h3f3c0315; // action70:  0.73442203
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3fe9b1ea; // action71:  1.82574201
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3f596a63; // action72:  0.84927958
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3ee84231; // action73:  0.45363000
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3f862983; // action74:  1.04814184
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3f891664; // action75:  1.07099581
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'hbe8a62bf; // action76: -0.27028462
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbf3ec1db; // action77: -0.74514550
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbf8bc5b1; // action78: -1.09197056
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbc7cbead; // action79: -0.01542632
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'hbe806bcf; // action80: -0.25082251
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3fb3c939; // action81:  1.40457833
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h3f17bd74; // action82:  0.59273458
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h3f83bcf0; // action83:  1.02920341
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbf7320c9; // action84: -0.94971901
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbfe023c1; // action85: -1.75109112
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'hbf89c961; // action86: -1.07645810
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3f58bb14; // action87:  0.84660459
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbfdb86db; // action88: -1.71505296
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbfaa5869; // action89: -1.33082306
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3f03579b; // action90:  0.51305550
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3faab5f5; // action91:  1.33367789
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbf27c1d5; // action92: -0.65530139
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'hbf8265f8; // action93: -1.01873684
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3efcb343; // action94:  0.49355516
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'hbf343345; // action95: -0.70390731
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'hbfd431f7; // action96: -1.65777481
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3edd787a; // action97:  0.43255979
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbd837e6d; // action98: -0.06420598
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3fd7e8a0; // action99:  1.68678665
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'hbed073a3; // action100: -0.40713224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h3fe9f7a9; // action101:  1.82787049
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'hbf52fa18; // action102: -0.82412863
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbf4175b4; // action103: -0.75570226
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h3ff1c003; // action104:  1.88867223
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbf5b3b25; // action105: -0.85637122
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3f343c0e; // action106:  0.70404136
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbf47cc67; // action107: -0.78046268
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'hbb0757a3; // action108: -0.00206516
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3fdc781a; // action109:  1.72241521
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'hbfbd8b11; // action110: -1.48080647
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h3fd88739; // action111:  1.69162667
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3fea0095; // action112:  1.82814276
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h3ff33027; // action113:  1.89990699
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'hbfc5c8ae; // action114: -1.54518676
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3fe85df6; // action115:  1.81536746
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3f0064de; // action116:  0.50153911
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3f07cbc1; // action117:  0.53045279
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3f6904fd; // action118:  0.91023237
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3f254b08; // action119:  0.64567614
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h3eefb0a1; // action120:  0.46814445
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3e9d6129; // action121:  0.30738190
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h3fe6968a; // action122:  1.80146909
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3ffb5d57; // action123:  1.96378601
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'hbf883440; // action124: -1.06409454
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'hbed717d9; // action125: -0.42010382
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h3f93b9f0; // action126:  1.15411186
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'hbfa8d3cb; // action127: -1.31896341
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h3f15cea5; // action128:  0.58518440
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3f3c45af; // action129:  0.73543829
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h3ec14554; // action130:  0.37748206
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbed2e11e; // action131: -0.41187376
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h3ee5f1ce; // action132:  0.44911045
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3cf7199d; // action133:  0.03016358
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'hbe91ee20; // action134: -0.28501987
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h3da14504; // action135:  0.07874492
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h3f592251; // action136:  0.84817988
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h3fa1f882; // action137:  1.26539636
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h3f3c59a8; // action138:  0.73574305
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h3fe4edba; // action139:  1.78850484
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h3f958d2d; // action140:  1.16837084
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h3d250c26; // action141:  0.04029479
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'hbed530b1; // action142: -0.41638711
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h3e270f53; // action143:  0.16314439
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'hbf7bd233; // action144: -0.98367614
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'hbf9d299a; // action145: -1.22783208
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h3fa623da; // action146:  1.29796910
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h3fb1eb85; // action147:  1.38999999
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3e783d7a; // action148:  0.24242201
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbf20aa62; // action149: -0.62759984
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'hbfb1fb8f; // action150: -1.39048946
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h3f7670dd; // action151:  0.96265966
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3ec7d11b; // action152:  0.39026722
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3f44c010; // action153:  0.76855564
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'hbd75d16e; // action154: -0.06001418
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h3f35f78d; // action155:  0.71080858
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbf427862; // action156: -0.75964940
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbe01bf26; // action157: -0.12670574
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbfbab0c6; // action158: -1.45851970
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'hbf99acf9; // action159: -1.20059121
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h3fb3f5ed; // action160:  1.40594256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h3f360a37; // action161:  0.71109337
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'hbee38b7f; // action162: -0.44442365
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'hbfcc0b09; // action163: -1.59408677
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h3e9a3204; // action164:  0.30116284
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'hbf426e09; // action165: -0.75949150
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbfe6e489; // action166: -1.80384934
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbfd41a5f; // action167: -1.65705478
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3d21c8d0; // action168:  0.03949815
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbf16eb35; // action169: -0.58952647
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbf5b925e; // action170: -0.85770214
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3f813800; // action171:  1.00952148
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'hbf00a36b; // action172: -0.50249356
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'hbf5eedca; // action173: -0.87081587
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3f0424e6; // action174:  0.51618803
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'hbe9ad916; // action175: -0.30243748
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'hbfcc298e; // action176: -1.59501815
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h3fdb46bf; // action177:  1.71309650
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h3f9ef04a; // action178:  1.24170804
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h3ff29cd5; // action179:  1.89541113
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h3e9f02f8; // action180:  0.31056952
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbec14420; // action181: -0.37747288
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h3f92d84c; // action182:  1.14722586
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h3eec811a; // action183:  0.46192247
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'hbfc1f94e; // action184: -1.51542068
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbfb663dd; // action185: -1.42492259
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'hbf9c1927; // action186: -1.21951759
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h3fd56843; // action187:  1.66724432
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h3f847169; // action188:  1.03471100
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbfc24a73; // action189: -1.51789701
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'hbfccb0d9; // action190: -1.59914696
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h3f39ef96; // action191:  0.72631204

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 5:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbfe5c153; // action0: -1.79496229
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3e5c9743; // action1:  0.21542077
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'hbedc44a2; // action2: -0.43021113
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3e0981b2; // action3:  0.13428381
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3f52bb76; // action4:  0.82317293
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbfbee69f; // action5: -1.49141300
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'hbfe0a4ba; // action6: -1.75502706
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h3fd5b335; // action7:  1.66953146
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'hbe2ecbbf; // action8: -0.17069910
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbf0f9fe8; // action9: -0.56103373
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h3ee3a9e7; // action10:  0.44465563
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbf985941; // action11: -1.19022381
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h3f279c47; // action12:  0.65472835
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h3e0d173c; // action13:  0.13778394
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h3fcaa2e2; // action14:  1.58309579
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'hbee4328c; // action15: -0.44569814
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h3d0983a5; // action16:  0.03357281
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'hbec60df0; // action17: -0.38682508
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h3ffca6d6; // action18:  1.97384143
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbf480bc8; // action19: -0.78142977
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'hbe67b367; // action20: -0.22627030
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbfe272a6; // action21: -1.76912379
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h3f79d7ab; // action22:  0.97594708
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbcab818e; // action23: -0.02093580
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbece4abd; // action24: -0.40291396
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3fc305dd; // action25:  1.52361643
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h3f9de825; // action26:  1.23364699
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3f41f897; // action27:  0.75769943
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'hbf97207c; // action28: -1.18067884
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbfe2e083; // action29: -1.77247655
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3f61ad91; // action30:  0.88155466
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h3fc6d565; // action31:  1.55338728
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbf89eaae; // action32: -1.07747436
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'hbf6a0532; // action33: -0.91414177
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'hbe9ac2e1; // action34: -0.30226806
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3dc6fcd8; // action35:  0.09716195
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'hbf90e762; // action36: -1.13206124
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'hbf118070; // action37: -0.56836605
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbfef1f6f; // action38: -1.86814678
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h3fdea6b0; // action39:  1.73946190
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3f337c94; // action40:  0.70111966
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h3f5ef274; // action41:  0.87088704
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3fbed54e; // action42:  1.49088454
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h3eb3c498; // action43:  0.35110927
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3f35c16d; // action44:  0.70998269
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'hbfbeea7b; // action45: -1.49153078
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h3f7d49f3; // action46:  0.98940963
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3f827cd2; // action47:  1.01943421
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h3f951d0e; // action48:  1.16494918
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbff154d9; // action49: -1.88540184
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h3f727891; // action50:  0.94715220
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbf874c89; // action51: -1.05702317
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h3f1a076c; // action52:  0.60167575
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'hbfb8e55a; // action53: -1.44449925
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'hbff8d254; // action54: -1.94391870
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'hbffd60d9; // action55: -1.97951806
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h3ea782ee; // action56:  0.32717079
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbfb4645d; // action57: -1.40931284
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3e18adc7; // action58:  0.14910041
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'hbfe06683; // action59: -1.75312841
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h3f9e1005; // action60:  1.23486388
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3fbef5ef; // action61:  1.49188030
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3cc76c9b; // action62:  0.02434378
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3fd3f611; // action63:  1.65594685
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3dbfcbf7; // action64:  0.09365075
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'hbe8194ae; // action65: -0.25308746
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbfef8d34; // action66: -1.87149668
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h3f83e278; // action67:  1.03034878
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3f0c2986; // action68:  0.54750860
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3f2e467c; // action69:  0.68076301
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h3fe645b5; // action70:  1.79900229
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3f4380fc; // action71:  0.76368690
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3e9f5b80; // action72:  0.31124496
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'hbf8418e2; // action73: -1.03200936
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'hbffbe39d; // action74: -1.96788371
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3d83c780; // action75:  0.06434536
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h3fcc25de; // action76:  1.59490561
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbf27d3c6; // action77: -0.65557516
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h3e382e96; // action78:  0.17986521
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbffc487c; // action79: -1.97096205
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3f15de81; // action80:  0.58542639
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3ff3c947; // action81:  1.90458000
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h3fd0be24; // action82:  1.63080263
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'hbf9b1388; // action83: -1.21153355
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbce1e0f6; // action84: -0.02757309
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h3ff99dc5; // action85:  1.95012724
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'hbf589e92; // action86: -0.84616959
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'hbe8ca9e3; // action87: -0.27473363
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h3ea9d34e; // action88:  0.33169025
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h3fb9da65; // action89:  1.45197737
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3f8053bb; // action90:  1.00255525
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3f12409d; // action91:  0.57129842
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h3f97b3c6; // action92:  1.18517375
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h3f82a8fb; // action93:  1.02078187
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3edcff34; // action94:  0.43163455
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'hbe84785c; // action95: -0.25873077
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h3f969629; // action96:  1.17645752
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3e0aa2fc; // action97:  0.13538736
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbfd5a18c; // action98: -1.66899252
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'hbe02d31b; // action99: -0.12775843
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'hbf480f1c; // action100: -0.78148055
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'hbfcd0e83; // action101: -1.60200536
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3fae9b6d; // action102:  1.36411822
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbf472bf0; // action103: -0.77801418
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h3fe56270; // action104:  1.79206657
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h3f51aff8; // action105:  0.81909132
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'hbfd18bb0; // action106: -1.63707542
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbfdfe0ba; // action107: -1.74904561
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3d2c0a7a; // action108:  0.04200218
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3f7c4503; // action109:  0.98542804
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h3fefd888; // action110:  1.87379551
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbf935fb9; // action111: -1.15135872
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3fe13714; // action112:  1.75949335
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'hbfefec1d; // action113: -1.87439311
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'hbf2fa4eb; // action114: -0.68611020
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3ef683b6; // action115:  0.48147362
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3f6a576f; // action116:  0.91539663
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3fd4ecce; // action117:  1.66347671
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3e79625c; // action118:  0.24353927
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3fdc63af; // action119:  1.72179210
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'hbfa12d4f; // action120: -1.25919521
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'hbfe5cb13; // action121: -1.79525983
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h3effcb91; // action122:  0.49959996
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3e04d628; // action123:  0.12972319
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3ea98e3f; // action124:  0.33116338
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'hbdf5af2f; // action125: -0.11996304
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h3fc4e248; // action126:  1.53815556
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'hbf9f3066; // action127: -1.24366450
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h3d50e667; // action128:  0.05100098
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'hbfba70fd; // action129: -1.45657313
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h3f9bd120; // action130:  1.21731949
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbf921f6a; // action131: -1.14158368
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'hbeead86f; // action132: -0.45868251
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3f8b1be8; // action133:  1.08678913
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'hbf47615c; // action134: -0.77882934
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h3fd9c260; // action135:  1.70124435
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'hbfa48abb; // action136: -1.28548372
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h3fc93188; // action137:  1.57182407
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'hbfc538d8; // action138: -1.54079723
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h3f5521df; // action139:  0.83254808
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'hbefde6e4; // action140: -0.49590218
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h3f0af290; // action141:  0.54276371
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3ec495c4; // action142:  0.38395512
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h3f26bd7d; // action143:  0.65132886
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3f6e99b0; // action144:  0.93203259
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h3eb7a400; // action145:  0.35867310
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'hbe2a5585; // action146: -0.16634186
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbfb67b9c; // action147: -1.42564726
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3f1b9d66; // action148:  0.60787046
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbfd716a1; // action149: -1.68037808
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'hbf769e96; // action150: -0.96335733
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h3fc64263; // action151:  1.54890096
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3fed6627; // action152:  1.85467994
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'hbfbcf771; // action153: -1.47630131
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h3f8984fd; // action154:  1.07437098
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'hbec8e98b; // action155: -0.39240679
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h3f80d998; // action156:  1.00664043
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbf212747; // action157: -0.62950557
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbe0c3c06; // action158: -0.13694772
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'hbfacf858; // action159: -1.35132885
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h3eb18d19; // action160:  0.34677961
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h3f451869; // action161:  0.76990372
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h3f04a224; // action162:  0.51809907
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'hbfd19252; // action163: -1.63727784
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbf77a1fa; // action164: -0.96731532
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3fefd87b; // action165:  1.87379396
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbf838762; // action166: -1.02756906
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h3f4bbf24; // action167:  0.79588532
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'hbe8a5d5b; // action168: -0.27024350
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbcedf9d9; // action169: -0.02904980
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbf871c96; // action170: -1.05555987
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3f069454; // action171:  0.52570081
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3fee9583; // action172:  1.86393774
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3f5e1bd8; // action173:  0.86761236
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'hbfe80284; // action174: -1.81257677
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'hbf812f72; // action175: -1.00926042
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3f8d4747; // action176:  1.10373771
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h3ff17774; // action177:  1.88645792
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbf9b2c84; // action178: -1.21229601
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbeb76ccf; // action179: -0.35825202
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h3dd8ad5c; // action180:  0.10579941
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbdf8cb58; // action181: -0.12148160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbfcbf08a; // action182: -1.59327817
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'hbefba5d6; // action183: -0.49149960
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'hbf1d3beb; // action184: -0.61419553
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbdbba4c9; // action185: -0.09162290
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'hbdf4d103; // action186: -0.11953928
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'hbfe6155e; // action187: -1.79752707
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h3fe2e7bf; // action188:  1.77269733
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbea3a9ad; // action189: -0.31965390
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'hbfb22221; // action190: -1.39166653
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h3fa562ca; // action191:  1.29207730

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 6:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbf3857e5; // action0: -0.72009116
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3e736b8e; // action1:  0.23771498
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'hbfdd29ef; // action2: -1.72784221
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3f1da4ce; // action3:  0.61579597
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3ff5eea2; // action4:  1.92134500
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h3fe9bb11; // action5:  1.82602131
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'hbf5c4a13; // action6: -0.86050528
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbf4581e0; // action7: -0.77151299
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h3f0241a1; // action8:  0.50881392
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbf764003; // action9: -0.96191424
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'hbf54929a; // action10: -0.83036196
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h3f96f798; // action11:  1.17943096
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'hbfe8cb17; // action12: -1.81869781
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h3fbb0dc6; // action13:  1.46135783
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h3fed3956; // action14:  1.85331225
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'hbfd5e925; // action15: -1.67117751
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'hbfebad3f; // action16: -1.84122455
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'hbffeb8ed; // action17: -1.99001849
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h3f44a206; // action18:  0.76809728
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbfc48b94; // action19: -1.53550959
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'hbfeedd74; // action20: -1.86613321
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h3f5a9f62; // action21:  0.85399449
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'hbffbc093; // action22: -1.96681440
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h3d4f2752; // action23:  0.05057461
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbf3e9974; // action24: -0.74452901
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3cffab0b; // action25:  0.03120949
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h3efae492; // action26:  0.49002510
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3ffe93b8; // action27:  1.98888302
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3fb1e810; // action28:  1.38989449
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h3f7708d3; // action29:  0.96497840
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3e921d76; // action30:  0.28538102
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbddef071; // action31: -0.10885704
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbfcfb129; // action32: -1.62259400
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3f813dfd; // action33:  1.00970423
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h3fa15847; // action34:  1.26050651
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'hbe856749; // action35: -0.26055363
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3f662209; // action36:  0.89895684
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h3e773647; // action37:  0.24141799
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbfcc96ce; // action38: -1.59835219
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h3facae68; // action39:  1.34907246
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3fb6449d; // action40:  1.42396891
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbfd8dffa; // action41: -1.69433522
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'hbf95ce75; // action42: -1.17036307
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbfb0615d; // action43: -1.37797129
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'hbda16846; // action44: -0.07881217
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3f8b1f13; // action45:  1.08688581
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbf79ea1e; // action46: -0.97622859
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'hbff26736; // action47: -1.89377475
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h3dfeba3d; // action48:  0.12437866
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbf7e18e8; // action49: -0.99256754
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h3f8a1ac0; // action50:  1.07894135
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbf5919bf; // action51: -0.84804910
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbfb188cf; // action52: -1.38698757
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'hbf772328; // action53: -0.96538019
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3fa78f99; // action54:  1.30906975
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h3edfdefd; // action55:  0.43724814
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h3f976b1b; // action56:  1.18295610
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbff4fe44; // action57: -1.91400957
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3ed662a8; // action58:  0.41872144
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'hbf80caaf; // action59: -1.00618541
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbf873352; // action60: -1.05625367
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'hbfa81714; // action61: -1.31320429
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'hbf2137ce; // action62: -0.62975776
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3f2063c9; // action63:  0.62652260
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3f9232bd; // action64:  1.14217341
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3f20abc1; // action65:  0.62762076
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h3f2d5c0d; // action66:  0.67718583
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbf40e84d; // action67: -0.75354463
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3e9cafb6; // action68:  0.30602807
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3fd1cf36; // action69:  1.63913608
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h3f0e31e2; // action70:  0.55544865
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3f9c22f3; // action71:  1.21981657
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'hbfa54a0d; // action72: -1.29132235
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'hbfd0b404; // action73: -1.63049364
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3f85c713; // action74:  1.04513776
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3ecfa4d0; // action75:  0.40555429
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h3e4cd0c3; // action76:  0.20001511
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbfaff36d; // action77: -1.37461627
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbf2d575e; // action78: -0.67711437
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbf270498; // action79: -0.65241385
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3f0496d9; // action80:  0.51792675
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3f381993; // action81:  0.71914023
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h3fe4545d; // action82:  1.78382456
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h3eca9d56; // action83:  0.39573163
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h3e88e795; // action84:  0.26739183
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h3f76e77b; // action85:  0.96446961
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'hbd6a28de; // action86: -0.05716788
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'hbd2d9f73; // action87: -0.04238839
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h3e72f857; // action88:  0.23727547
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h3f50f0a4; // action89:  0.81617188
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3f840b77; // action90:  1.03159988
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3e97fe20; // action91:  0.29686069
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbee332ee; // action92: -0.44374794
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h3f9148c6; // action93:  1.13503337
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3f39b068; // action94:  0.72534800
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'hbf8db178; // action95: -1.10697842
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h3ed8b112; // action96:  0.42322594
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3fcdde3d; // action97:  1.60834467
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbfc1f1aa; // action98: -1.51518750
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3fb02755; // action99:  1.37620032
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h3fa01851; // action100:  1.25074208
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h3dd03cc7; // action101:  0.10167842
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3fc2bc0c; // action102:  1.52136374
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbfd473e8; // action103: -1.65978718
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'hbf813dae; // action104: -1.00969481
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbf2b29c4; // action105: -0.66860604
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3fdf7002; // action106:  1.74560571
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h3f838b68; // action107:  1.02769184
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3fd16fd9; // action108:  1.63622582
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3dc0ed83; // action109:  0.09420302
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'hbfffd447; // action110: -1.99866569
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h3f88cfca; // action111:  1.06884122
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'hbffa9913; // action112: -1.95779645
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'hbf80ae36; // action113: -1.00531650
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h3feff33a; // action114:  1.87461019
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3fd86125; // action115:  1.69046462
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3faec939; // action116:  1.36551583
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'hbf806c12; // action117: -1.00329804
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3f469a63; // action118:  0.77579325
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'hbd8c7f4a; // action119: -0.06860216
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'hbf9d9dfc; // action120: -1.23138380
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'hbfa34161; // action121: -1.27543271
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'hbfb74317; // action122: -1.43173492
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3fa61859; // action123:  1.29761803
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'hbf5f4da6; // action124: -0.87227857
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h3e5be289; // action125:  0.21473135
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbfe8588f; // action126: -1.81520259
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3f60a947; // action127:  0.87758297
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h3fd8a3be; // action128:  1.69249701
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3e9601fd; // action129:  0.29298392
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'hbf659d02; // action130: -0.89692700
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h3f85638d; // action131:  1.04210055
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h3f3d0d49; // action132:  0.73848397
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'hbf4451cc; // action133: -0.76687312
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3f141286; // action134:  0.57840765
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'hbffaf068; // action135: -1.96046162
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'hbfe38543; // action136: -1.77750432
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'hbff2c4c9; // action137: -1.89663041
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h3fc92059; // action138:  1.57129967
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'hbfc01f6e; // action139: -1.50095916
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'hbfb88a59; // action140: -1.44172204
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'hbfc3569c; // action141: -1.52608061
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'hbfd8f935; // action142: -1.69510520
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h3eebaec4; // action143:  0.46031773
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3ee5ee87; // action144:  0.44908544
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h3f213e60; // action145:  0.62985802
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'hbf34a4ef; // action146: -0.70564169
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h3fa65d22; // action147:  1.29971719
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'hbf12b810; // action148: -0.57312107
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h3f2fbf26; // action149:  0.68651044
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h3f3134a7; // action150:  0.69220966
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbf983f7d; // action151: -1.18943751
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3e085944; // action152:  0.13315302
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3f8a5fe8; // action153:  1.08105183
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h3ffade26; // action154:  1.95990443
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h3fa67e44; // action155:  1.30072832
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbfe04d4b; // action156: -1.75235879
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbeff98b7; // action157: -0.49921200
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbfaee1d0; // action158: -1.36626625
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'hbfb5d283; // action159: -1.42048681
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbfdfcc8c; // action160: -1.74842978
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h3f5cbc08; // action161:  0.86224413
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'hbf9af0ac; // action162: -1.21046972
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'hbe8ad93c; // action163: -0.27118862
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbeeb005b; // action164: -0.45898709
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3db4c923; // action165:  0.08827426
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h3fd0c442; // action166:  1.63098931
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbfa15cac; // action167: -1.26064062
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3ec415df; // action168:  0.38297936
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h3fffaa8a; // action169:  1.99739194
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbf97ee4a; // action170: -1.18695951
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3fdde65d; // action171:  1.73359263
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3fd681aa; // action172:  1.67583203
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3fbda6c7; // action173:  1.48165214
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3e4eab8d; // action174:  0.20182629
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3ec02af1; // action175:  0.37532762
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3f9863ba; // action176:  1.19054341
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h3f8ff9e1; // action177:  1.12481320
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h3e2b14bb; // action178:  0.16707127
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbff86421; // action179: -1.94055569
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'hbfd9c985; // action180: -1.70146239
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbfebd8d9; // action181: -1.84255517
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbfc2f848; // action182: -1.52320194
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'hbf0ea6a2; // action183: -0.55723011
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3fcfa85b; // action184:  1.62232530
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbff8f9e7; // action185: -1.94512641
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3f57ddb3; // action186:  0.84322661
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h3ff3d65a; // action187:  1.90497899
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbfbc91bb; // action188: -1.47319734
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbfde1b59; // action189: -1.73520958
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h3f8c423e; // action190:  1.09577155
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'hbf3ef567; // action191: -0.74593204

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 7:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbfac2ebe; // action0: -1.34517646
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3fcfef13; // action1:  1.62448347
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3fc19bab; // action2:  1.51256311
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3df56564; // action3:  0.11982229
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3fc48da4; // action4:  1.53557253
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h3e870607; // action5:  0.26371786
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3ed82845; // action6:  0.42218223
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbfc4af6c; // action7: -1.53660345
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h3e0600dd; // action8:  0.13086267
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbf1e82f5; // action9: -0.61918575
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h3e7d2c61; // action10:  0.24723960
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbee4f624; // action11: -0.44719040
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'hbf08eff7; // action12: -0.53491157
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbfc93cdb; // action13: -1.57216966
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbfc21224; // action14: -1.51617861
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3f5f4ef6; // action15:  0.87229860
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h3fe6621d; // action16:  1.79986918
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h3f4253a0; // action17:  0.75908852
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h3f4d26bf; // action18:  0.80137247
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbf4ef35f; // action19: -0.80840105
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h3f7148ec; // action20:  0.94251895
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h3fd40593; // action21:  1.65642011
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h3fa8a633; // action22:  1.31757200
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h3edf1acc; // action23:  0.43575132
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h3f842702; // action24:  1.03244042
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3fe1b389; // action25:  1.76329148
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'hbf145dd2; // action26: -0.57955658
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'hbfea305d; // action27: -1.82960093
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'hbf8f7570; // action28: -1.12077141
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbfa65820; // action29: -1.29956436
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'hbfc7ca8f; // action30: -1.56086910
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h3ff8c2ee; // action31:  1.94344878
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbfa52646; // action32: -1.29023051
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3fa3e2d0; // action33:  1.28035927
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h3fc77be3; // action34:  1.55846822
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3f5e65cb; // action35:  0.86874074
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'hbf87c336; // action36: -1.06064487
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'hbf22f340; // action37: -0.63652420
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbfdad61c; // action38: -1.70965910
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h3f6760f6; // action39:  0.90382326
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3f6c250c; // action40:  0.92244029
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbffdee73; // action41: -1.98383939
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3fcb9c02; // action42:  1.59069848
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h3f8f58a0; // action43:  1.11989212
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'hbe11fbed; // action44: -0.14256258
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3e070944; // action45:  0.13187128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbfaa8fa8; // action46: -1.33250904
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'hbff40279; // action47: -1.90632546
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h3fa5dbed; // action48:  1.29577410
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbee8b67e; // action49: -0.45451730
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbfce6e5f; // action50: -1.61274326
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbf2fbed4; // action51: -0.68650556
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbf23c7de; // action52: -0.63976848
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'hbf732ed0; // action53: -0.94993305
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3e324452; // action54:  0.17408875
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h3fa9393e; // action55:  1.32205939
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h3ffa6765; // action56:  1.95628035
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbe769538; // action57: -0.24080360
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'hbe7e43d5; // action58: -0.24830563
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'hbda3ade9; // action59: -0.07992155
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbfade6b7; // action60: -1.35860336
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3fc23ef5; // action61:  1.51754630
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3fe08276; // action62:  1.75398135
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3fc26741; // action63:  1.51877606
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'hbfe857d6; // action64: -1.81518054
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3ee45c9d; // action65:  0.44601908
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbe12dec3; // action66: -0.14342789
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h3fe8cdbe; // action67:  1.81877875
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3ff5e1cc; // action68:  1.92095327
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3fa39719; // action69:  1.27804863
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'hbf37f062; // action70: -0.71851170
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'hbe6dd4ca; // action71: -0.23225704
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3f9eb7ad; // action72:  1.23998034
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'hbd7df849; // action73: -0.06200436
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3f9986a8; // action74:  1.19942188
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'hbf26f4dc; // action75: -0.65217376
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h3fbedf8d; // action76:  1.49119723
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbf7f9367; // action77: -0.99834293
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbf06cdf5; // action78: -0.52658015
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbf4ddf54; // action79: -0.80418897
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'hbfd80890; // action80: -1.68776131
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'hbdb0e314; // action81: -0.08637062
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'hbfae3d2a; // action82: -1.36124158
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'hbffd3cdc; // action83: -1.97841978
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbf0d7a38; // action84: -0.55264616
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h3f7fd091; // action85:  0.99927622
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h3e93429a; // action86:  0.28761750
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3fe297e1; // action87:  1.77025998
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h3f04403d; // action88:  0.51660520
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbfc73e37; // action89: -1.55658615
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'hbf64ca51; // action90: -0.89371210
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'hbf95b80c; // action91: -1.16967916
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h3ecb361b; // action92:  0.39689717
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h3fb40e46; // action93:  1.40668559
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'hbe4faa51; // action94: -0.20279814
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h3f95c664; // action95:  1.17011690
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'hbff928ea; // action96: -1.94656110
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'hbfada548; // action97: -1.35660648
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbf0f2e4f; // action98: -0.55930036
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3fbefe89; // action99:  1.49214280
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h3f5d99f8; // action100:  0.86563063
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'hbf92ca59; // action101: -1.14680016
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3f7cd3e6; // action102:  0.98760831
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbf82563e; // action103: -1.01825690
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'hbfd63e37; // action104: -1.67377365
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbff95db1; // action105: -1.94817173
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'hbc369197; // action106: -0.01114311
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbfcc61e1; // action107: -1.59673703
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3edc2b27; // action108:  0.43001673
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3d26b8dc; // action109:  0.04070364
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h3fd604e5; // action110:  1.67202437
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h3ecf72e6; // action111:  0.40517348
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'hbf8b364a; // action112: -1.08759427
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h3fe8b098; // action113:  1.81788921
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h3f0a8f3e; // action114:  0.54124820
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'hbf06df54; // action115: -0.52684522
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'hbfd26fcd; // action116: -1.64403689
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3f6fae4c; // action117:  0.93625331
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'hbfa13e92; // action118: -1.25972199
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'hbfdba884; // action119: -1.71608019
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h3fa80d93; // action120:  1.31291425
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3fa9880f; // action121:  1.32446468
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'hbe303277; // action122: -0.17206751
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3f96a877; // action123:  1.17701614
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3fd84c31; // action124:  1.68982518
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'hbfc1a6c7; // action125: -1.51290214
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbf79e97a; // action126: -0.97621882
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3fdc7100; // action127:  1.72219849
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h3f220011; // action128:  0.63281351
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3f0c1411; // action129:  0.54718119
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'hbf4ef88b; // action130: -0.80847996
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbfe492ae; // action131: -1.78572631
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h3f77c35d; // action132:  0.96782476
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3fdef4bf; // action133:  1.74184406
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3eb1e26e; // action134:  0.34743065
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h3e7d5984; // action135:  0.24741179
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'hbf5b6330; // action136: -0.85698223
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h3f57b6b1; // action137:  0.84263140
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'hbf542841; // action138: -0.82873923
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'hbea2c33f; // action139: -0.31789586
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h3f8c90e0; // action140:  1.09817123
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h3fc69494; // action141:  1.55140924
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3f9e287e; // action142:  1.23561072
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h3fb57560; // action143:  1.41764450
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3f92e0ed; // action144:  1.14748919
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h3fbb6974; // action145:  1.46415567
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h3e363fce; // action146:  0.17797777
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h3ee195b3; // action147:  0.44059524
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3f1c28c0; // action148:  0.60999680
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbef330ed; // action149: -0.47498265
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h3fdba84d; // action150:  1.71607363
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h3f98971d; // action151:  1.19211161
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3f19780a; // action152:  0.59948790
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3fbf4825; // action153:  1.49438918
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h3f060953; // action154:  0.52357978
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'hbfd3bd58; // action155: -1.65421581
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h3fbc9a7c; // action156:  1.47346449
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h3fc84720; // action157:  1.56467056
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h3f8b3688; // action158:  1.08760166
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'hbfeec1cf; // action159: -1.86528957
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbfccb472; // action160: -1.59925675
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'hbf14be87; // action161: -0.58103222
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h3fa31846; // action162:  1.27417827
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'hbfc86030; // action163: -1.56543541
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbf945409; // action164: -1.15881455
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3fcf9b88; // action165:  1.62193394
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbf39f4c4; // action166: -0.72639108
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbf8f6322; // action167: -1.12021279
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3fcdba7d; // action168:  1.60725367
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbea5cffc; // action169: -0.32385242
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbfe171be; // action170: -1.76128364
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3fc770be; // action171:  1.55812812
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3f7dc9f9; // action172:  0.99136311
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'hbfb3c5ba; // action173: -1.40447164
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3f547fc9; // action174:  0.83007485
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'hbfe90110; // action175: -1.82034492
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'hbe958273; // action176: -0.29201087
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'hbf37c9fa; // action177: -0.71792567
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h3ea1dd95; // action178:  0.31614366
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbf8a891d; // action179: -1.08230937
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'hbf12c526; // action180: -0.57332075
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h3fc2d2f4; // action181:  1.52206278
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbff37030; // action182: -1.90186119
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h3f26b3e3; // action183:  0.65118235
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3e96c062; // action184:  0.29443651
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbefafd73; // action185: -0.49021491
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'hbf9d413e; // action186: -1.22855353
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'hbdbe6cff; // action187: -0.09298133
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h3f92b3c3; // action188:  1.14611089
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbfad19d5; // action189: -1.35235083
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h3fafb72e; // action190:  1.37277770
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'hbf43a7b2; // action191: -0.76427758

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 8:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbfe23f9c; // action0: -1.76756620
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'hbf941c9c; // action1: -1.15712309
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'hbf0856eb; // action2: -0.53257626
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'hbfdadd73; // action3: -1.70988309
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'hbf76582b; // action4: -0.96228284
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h3fb086a7; // action5:  1.37910926
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3e913bdd; // action6:  0.28365985
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbf2b8e43; // action7: -0.67013949
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'hbea5eefd; // action8: -0.32408896
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbf98e401; // action9: -1.19445813
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h3c5ebf69; // action10:  0.01359544
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h3fa4e5ad; // action11:  1.28825915
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'hbf8b6a2d; // action12: -1.08917773
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h3f613871; // action13:  0.87976748
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h3f2fbf7f; // action14:  0.68651575
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'hbff45858; // action15: -1.90894604
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'hbdeb53d8; // action16: -0.11490601
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'hbf1db844; // action17: -0.61609292
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'hbfa0ad3c; // action18: -1.25528669
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h3f141c12; // action19:  0.57855332
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'hbdcb8f14; // action20: -0.09939399
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h3f927469; // action21:  1.14417756
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'hbfbb7af2; // action22: -1.46468949
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbed61252; // action23: -0.41810852
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbfa252c2; // action24: -1.26815057
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3f2f8ab7; // action25:  0.68571037
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'hbfc89eed; // action26: -1.56735003
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'hbec755e6; // action27: -0.38932723
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'hbd31628b; // action28: -0.04330687
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbf598ac7; // action29: -0.84977382
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3f75566c; // action30:  0.95834994
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbfde5291; // action31: -1.73689473
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbfd1a96b; // action32: -1.63798273
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3ea5180e; // action33:  0.32244915
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h3fe93c1e; // action34:  1.82214713
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3faa7731; // action35:  1.33176243
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3f05116e; // action36:  0.51979721
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'hbfbc6613; // action37: -1.47186506
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbfad5652; // action38: -1.35419679
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'hbf52b51c; // action39: -0.82307601
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'hbfd3d4a0; // action40: -1.65492630
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h3fffb9ba; // action41:  1.99785542
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3fbff256; // action42:  1.49958301
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h3e87b7f5; // action43:  0.26507536
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3f91631a; // action44:  1.13583684
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'hbf3c4ba6; // action45: -0.73552930
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbe06b70d; // action46: -0.13155766
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3ff68854; // action47:  1.92603540
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h3e20b779; // action48:  0.15694989
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbefa3649; // action49: -0.48869541
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbfe7b859; // action50: -1.81031334
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h3ebd298a; // action51:  0.36945754
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbff2a3a0; // action52: -1.89561844
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h3f704f16; // action53:  0.93870676
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'hbfa15ee0; // action54: -1.26070786
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h3eb3dde1; // action55:  0.35130218
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h3f240925; // action56:  0.64076453
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbefd067b; // action57: -0.49419007
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'hbfce0e91; // action58: -1.60981953
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'hbfac52a0; // action59: -1.34627151
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbfa0291d; // action60: -1.25125468
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3e87794e; // action61:  0.26459736
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3f800b9d; // action62:  1.00035441
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3f85ffff; // action63:  1.04687488
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3f9acf98; // action64:  1.20946026
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3ecc5466; // action65:  0.39908141
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h3eff0320; // action66:  0.49807072
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h3fee1ea5; // action67:  1.86031020
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3f9c823c; // action68:  1.22272444
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'hbd31638a; // action69: -0.04330782
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'hbeeada62; // action70: -0.45869738
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'hbfd717d4; // action71: -1.68041468
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'hbf3a3bc1; // action72: -0.72747427
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'hbe80ac11; // action73: -0.25131276
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3ec839dc; // action74:  0.39106643
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3f7c4cc9; // action75:  0.98554665
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'hbf48bd2b; // action76: -0.78413647
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbfb14b8c; // action77: -1.38511801
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h3fd75d71; // action78:  1.68253911
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h3f46ec10; // action79:  0.77703953
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3f9fb46c; // action80:  1.24769354
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3dd3d42c; // action81:  0.10343203
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'hbffb8919; // action82: -1.96512139
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h3d9a7fac; // action83:  0.07543883
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h3f70eadd; // action84:  0.94108373
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h3fa8f9d4; // action85:  1.32012415
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h3ffa7f43; // action86:  1.95700872
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3dffbcbf; // action87:  0.12487172
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbfb537b7; // action88: -1.41576278
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbe04bf7b; // action89: -0.12963669
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3daf9e65; // action90:  0.08575133
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'hbff00771; // action91: -1.87522709
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbf2ac7ca; // action92: -0.66711104
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'hbfb4ed4a; // action93: -1.41349149
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3f803362; // action94:  1.00156808
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h3f8befce; // action95:  1.09325576
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h3fa6b611; // action96:  1.30243123
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3f65a5ce; // action97:  0.89706123
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h3fcccf04; // action98:  1.60006762
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3ebfa861; // action99:  0.37433150
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h3fbc67b0; // action100:  1.47191429
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'hbf14ee1d; // action101: -0.58175832
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'hbfc71980; // action102: -1.55546570
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h3fd3ff4e; // action103:  1.65622878
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'hbfcd275b; // action104: -1.60276353
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h3fa15673; // action105:  1.26045072
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'hbeaa2d29; // action106: -0.33237579
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h3f907db4; // action107:  1.12883615
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'hbff88787; // action108: -1.94163597
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3f8ca07b; // action109:  1.09864748
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'hbf83ba71; // action110: -1.02912724
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h3fd24b1f; // action111:  1.64291751
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'hbf001609; // action112: -0.50033623
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h3f739cbd; // action113:  0.95161039
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h3ef83430; // action114:  0.48477316
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3ffb3a09; // action115:  1.96270859
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3e81d9e1; // action116:  0.25361541
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'hbfc04bdc; // action117: -1.50231504
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3f8934fd; // action118:  1.07192957
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3e204013; // action119:  0.15649442
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'hbf721979; // action120: -0.94570118
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3f77ce6e; // action121:  0.96799362
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h3f64dece; // action122:  0.89402473
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'hbfc559fa; // action123: -1.54180837
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3ea1c21e; // action124:  0.31593412
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h3f8f035c; // action125:  1.11729002
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbf61ffa1; // action126: -0.88280684
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3ef7890e; // action127:  0.48346752
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h3f614475; // action128:  0.87995082
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3ffe0266; // action129:  1.98444819
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'hbfc55ff0; // action130: -1.54199028
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h3f8ff5d3; // action131:  1.12468946
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h3d5970fa; // action132:  0.05308626
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3cb6a599; // action133:  0.02229576
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'hbf71b694; // action134: -0.94419217
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'hbfb8b641; // action135: -1.44306195
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h3f37b5d4; // action136:  0.71761823
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'hbfcd9d00; // action137: -1.60635376
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'hbf88bc91; // action138: -1.06825459
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h3f21789a; // action139:  0.63074648
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h3fc3ad29; // action140:  1.52872193
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'hbfb78474; // action141: -1.43372965
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3feedcb3; // action142:  1.86611021
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'hbf3620db; // action143: -0.71143883
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3eb29584; // action144:  0.34879696
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h3ffc4d44; // action145:  1.97110796
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'hbf997e4d; // action146: -1.19916689
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbf3734be; // action147: -0.71564853
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3ff7c45f; // action148:  1.93568027
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbff629dd; // action149: -1.92315257
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h3ebcbee6; // action150:  0.36864394
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h3f29a3ec; // action151:  0.66265750
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'hbff66575; // action152: -1.92497122
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3fa16335; // action153:  1.26084006
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'hbf966c69; // action154: -1.17518342
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'hbf36e753; // action155: -0.71446723
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbfede5a8; // action156: -1.85857105
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h3fdb63c3; // action157:  1.71398199
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h3e46c393; // action158:  0.19410543
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'hbe71aa15; // action159: -0.23600037
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h3ea79a0a; // action160:  0.32734710
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h3f6454f4; // action161:  0.89192128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'hbfcf51cf; // action162: -1.61968410
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'hbfebc047; // action163: -1.84180534
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbfa8a51d; // action164: -1.31753886
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'hbf659eba; // action165: -0.89695323
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h3fdb05d2; // action166:  1.71111512
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbf712803; // action167: -0.94201678
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'hbe952e5e; // action168: -0.29136938
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h3f9a87b7; // action169:  1.20726669
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbfd12d89; // action170: -1.63420212
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'hbf98ce52; // action171: -1.19379640
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'hbfcc6a8e; // action172: -1.59700179
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3f9b4618; // action173:  1.21307659
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'hbfa2030a; // action174: -1.26571774
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'hbe805081; // action175: -0.25061420
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'hbf6f0aa4; // action176: -0.93375611
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h3fca093d; // action177:  1.57840693
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbfc533e0; // action178: -1.54064560
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbf1bf05c; // action179: -0.60913634
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h3f63f620; // action180:  0.89047432
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h3f8f2f9d; // action181:  1.11864054
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h3e68cb32; // action182:  0.22733763
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'hbfd18c1b; // action183: -1.63708818
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3fa944fc; // action184:  1.32241774
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h3ffca33f; // action185:  1.97373188
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3f121705; // action186:  0.57066375
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'hbf64674d; // action187: -0.89220124
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbff37fdd; // action188: -1.90233958
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbfa59b5e; // action189: -1.29380393
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h3f8cb55e; // action190:  1.09928489
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'hbe4f4775; // action191: -0.20242102

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 9:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbff6a522; // action0: -1.92691445
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3fddb0cf; // action1:  1.73195827
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3fde8646; // action2:  1.73847270
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'hbf8295f3; // action3: -1.02020109
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3f5baa01; // action4:  0.85806280
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbf8e5f45; // action5: -1.11228240
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3e11a557; // action6:  0.14223228
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h3f996b86; // action7:  1.19859385
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h3fd7ce1a; // action8:  1.68597722
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h3fb53257; // action9:  1.41559875
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'hbf0e1b9c; // action10: -0.55510879
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbf2db319; // action11: -0.67851406
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h3fa170f3; // action12:  1.26125944
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbe2b04bf; // action13: -0.16701029
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbfebdf75; // action14: -1.84275687
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'hbf80cb2c; // action15: -1.00620031
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'hbff265b3; // action16: -1.89372861
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'hbf85cd3d; // action17: -1.04532588
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h3f923ae1; // action18:  1.14242184
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbf11fe9e; // action19: -0.57029140
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h3f999c53; // action20:  1.20008314
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbe3f23f8; // action21: -0.18666065
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h3fb29ccd; // action22:  1.39541018
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbd3b812d; // action23: -0.04577749
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbdcfbe55; // action24: -0.10143725
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3fee7c6a; // action25:  1.86317182
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'hbf824777; // action26: -1.01780593
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'hbcf45ac0; // action27: -0.02982843
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'hbfe1e39e; // action28: -1.76475883
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbfd5db44; // action29: -1.67075396
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3fdcb4f1; // action30:  1.72427189
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbff8e4bc; // action31: -1.94448042
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbf5a632a; // action32: -0.85307562
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3fd9b846; // action33:  1.70093608
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h3fed3942; // action34:  1.85330987
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'hbf84640b; // action35: -1.03430307
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3e5fab10; // action36:  0.21842599
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'hbfd95fbf; // action37: -1.69823444
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbf973564; // action38: -1.18131685
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'hbeb65259; // action39: -0.35609701
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3de15df4; // action40:  0.11004248
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbfcaf94a; // action41: -1.58573270
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3f2a8a44; // action42:  0.66617227
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h3f8449fb; // action43:  1.03350770
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3f823e5e; // action44:  1.01752830
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'hbf8243b0; // action45: -1.01769066
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h3f56e166; // action46:  0.83937681
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'hbf7fae07; // action47: -0.99874920
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h3eea4d5b; // action48:  0.45762143
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbea29a57; // action49: -0.31758377
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h3e49daff; // action50:  0.19712447
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbff1a019; // action51: -1.88769829
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbfa5b569; // action52: -1.29459870
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h3fe976ab; // action53:  1.82393396
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3f3448eb; // action54:  0.70423764
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'hbeefcb6c; // action55: -0.46834886
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'hbf72f379; // action56: -0.94902760
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbfa5decf; // action57: -1.29586208
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'hbd15ec89; // action58: -0.03660253
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h3fe6c4ec; // action59:  1.80288458
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h3f124e0a; // action60:  0.57150328
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3fa23b0c; // action61:  1.26742697
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3f678ee8; // action62:  0.90452433
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3fefd9ac; // action63:  1.87383032
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3fb8f715; // action64:  1.44504035
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3fe02df2; // action65:  1.75140214
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbf9cc619; // action66: -1.22479546
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbfc6ded2; // action67: -1.55367494
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3f58daef; // action68:  0.84709066
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3fe1616e; // action69:  1.76078582
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h3b6bb093; // action70:  0.00359634
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3f67e697; // action71:  0.90586227
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'hbf04ba25; // action72: -0.51846534
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3fd2ec11; // action73:  1.64782917
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'hbf3dade4; // action74: -0.74093461
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'hbf11e527; // action75: -0.56990284
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'hbfa834bf; // action76: -1.31410968
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbfc64ca0; // action77: -1.54921341
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbfb06be0; // action78: -1.37829208
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbf986199; // action79: -1.19047844
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3f8c0583; // action80:  1.09391820
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3e87ade6; // action81:  0.26499861
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'hbed1f726; // action82: -0.41008872
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h3fb460ba; // action83:  1.40920186
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbfe9ed9f; // action84: -1.82756412
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h3ff35c94; // action85:  1.90126276
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h3e6d57bf; // action86:  0.23178004
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3f1d2727; // action87:  0.61387867
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbf4a2726; // action88: -0.78965986
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h3e899e4d; // action89:  0.26878586
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3f9ff6f9; // action90:  1.24972451
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3fd1ff54; // action91:  1.64060450
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbf85606c; // action92: -1.04200506
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h3f63d017; // action93:  0.88989395
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3d68a2c9; // action94:  0.05679587
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h3f15ebb8; // action95:  0.58562803
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'hbf71e031; // action96: -0.94482714
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3f7dc822; // action97:  0.99133503
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbfd2c49a; // action98: -1.64662480
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3f77c789; // action99:  0.96788841
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h3fc53102; // action100:  1.54055810
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h3f703b76; // action101:  0.93840730
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3fa30852; // action102:  1.27369142
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbd05bdd5; // action103: -0.03265174
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h3f922b62; // action104:  1.14194894
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbcc701d2; // action105: -0.02429286
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'hbfef0810; // action106: -1.86743355
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbfec427e; // action107: -1.84577918
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'hbfdc651e; // action108: -1.72183585
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3f0ad3a9; // action109:  0.54229218
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'hbec45aa1; // action110: -0.38350394
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbf0c035f; // action111: -0.54692644
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3fb1b861; // action112:  1.38843930
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h3f4b07f9; // action113:  0.79309040
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'hbfb51cd3; // action114: -1.41494215
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'hbf5b121b; // action115: -0.85574502
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'hbfc3128b; // action116: -1.52400339
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3fbeee16; // action117:  1.49164081
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'hbf1c4091; // action118: -0.61036021
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'hbf024e62; // action119: -0.50900853
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'hbeb59636; // action120: -0.35466164
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3e7371f2; // action121:  0.23773935
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h3fd41da5; // action122:  1.65715468
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3f9425a9; // action123:  1.15739930
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'hbf32668b; // action124: -0.69687718
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h3fce3fd7; // action125:  1.61132324
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbf84ec8e; // action126: -1.03846908
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'hbfd34715; // action127: -1.65060675
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'hbf82a362; // action128: -1.02061105
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'hbff9bfec; // action129: -1.95116949
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'hbfa82298; // action130: -1.31355572
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbfecbdd9; // action131: -1.84954369
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'hbfd23f2f; // action132: -1.64255321
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3e30253a; // action133:  0.17201701
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3f13aa9e; // action134:  0.57682216
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h3fff315b; // action135:  1.99369371
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h3feb96a4; // action136:  1.84053469
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'hbe59f53e; // action137: -0.21284959
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h3eb354d8; // action138:  0.35025668
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'hbfde2d2e; // action139: -1.73575377
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h3f6bc2b9; // action140:  0.92093998
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h3f2a8ba1; // action141:  0.66619307
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3f8ea513; // action142:  1.11441267
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h3fe1bda0; // action143:  1.76359940
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3cc19404; // action144:  0.02363015
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h3ea7b5ef; // action145:  0.32755992
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h3c3de8cf; // action146:  0.01159115
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h3f95b808; // action147:  1.16967869
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3edd22df; // action148:  0.43190667
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbf93b227; // action149: -1.15387428
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'hbf34681e; // action150: -0.70471370
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbf86d15d; // action151: -1.05326426
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3ec580b5; // action152:  0.38574758
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3cc15cc7; // action153:  0.02360381
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'hbfea7b4e; // action154: -1.83188796
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'hbf916adf; // action155: -1.13607395
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbfca9697; // action156: -1.58272064
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbea86cad; // action157: -0.32895413
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbf295064; // action158: -0.66138291
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h3f51c40e; // action159:  0.81939781
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbf8f3e9a; // action160: -1.11909795
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h3ed2762b; // action161:  0.41105780
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h3d7e9547; // action162:  0.06215408
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h3f91b761; // action163:  1.13840878
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbf9c2bb5; // action164: -1.22008383
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'hbfc6a333; // action165: -1.55185544
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h3f8997c2; // action166:  1.07494378
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h3f49e20e; // action167:  0.78860557
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3f5a790f; // action168:  0.85340971
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h3e235e29; // action169:  0.15953888
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h3fec4c5c; // action170:  1.84608030
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3ff91c1c; // action171:  1.94617033
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3fd5241b; // action172:  1.66516435
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3ef2255d; // action173:  0.47294131
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3f88ab5e; // action174:  1.06772971
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'hbf8d00fc; // action175: -1.10159254
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'hbe5ae260; // action176: -0.21375418
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'hbfa51343; // action177: -1.28965032
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbf896740; // action178: -1.07346344
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbe9e09ac; // action179: -0.30866754
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h3fa2ac1a; // action180:  1.27087712
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbe8b8098; // action181: -0.27246547
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h3dd3d2f6; // action182:  0.10342972
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'hbdf7a550; // action183: -0.12092078
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'hbf67486b; // action184: -0.90344876
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h3e9a167d; // action185:  0.30095282
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3f0bf5a4; // action186:  0.54671693
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'hbfda0024; // action187: -1.70312929
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbfef7f4c; // action188: -1.87107229
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h3e37fea9; // action189:  0.17968239
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h3fcbdaec; // action190:  1.59261847
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'hbfa9e6de; // action191: -1.32735801

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 10:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h3edb0842; // action0:  0.42779738
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'hbfbf1e2b; // action1: -1.49310815
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3f50017d; // action2:  0.81252271
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'hbfa2ed00; // action3: -1.27285767
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'hbfc77838; // action4: -1.55835629
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbf4cf9f1; // action5: -0.80068880
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'hbea88b88; // action6: -0.32918954
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h3e9ef1fb; // action7:  0.31043991
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'hbfa86539; // action8: -1.31558907
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h3ffff9c9; // action9:  1.99981034
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h3ff10aaf; // action10:  1.88313854
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbf6ddb39; // action11: -0.92912632
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'hbfd42c60; // action12: -1.65760422
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h3fe3ecbb; // action13:  1.78066194
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbfe9823b; // action14: -1.82428682
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3e9fed67; // action15:  0.31235811
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'hbf6cc771; // action16: -0.92491823
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'hbf96167d; // action17: -1.17256129
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h3e4a966e; // action18:  0.19783947
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbf6a4e15; // action19: -0.91525394
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h3f2ac708; // action20:  0.66709948
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbf820b4a; // action21: -1.01596951
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'hbf4286b1; // action22: -0.75986773
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbf18969d; // action23: -0.59604818
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h3fe89a11; // action24:  1.81720173
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3fa79424; // action25:  1.30920839
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h3f9ea804; // action26:  1.23950243
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3e5c09ec; // action27:  0.21488160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'hbf05827f; // action28: -0.52152246
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbe1b6efb; // action29: -0.15179054
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3efdd05b; // action30:  0.49573025
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h3ec6941a; // action31:  0.38784868
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbfe99aa8; // action32: -1.82503223
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3fc7e400; // action33:  1.56164551
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'hbfb2e984; // action34: -1.39775133
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'hbfe45827; // action35: -1.78394020
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3f8c9094; // action36:  1.09816217
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h3e858450; // action37:  0.26077509
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h3fa803c5; // action38:  1.31261504
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h3fe3292b; // action39:  1.77469385
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'hbfefd55b; // action40: -1.87369859
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h3d2f21be; // action41:  0.04275679
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'hbeed1858; // action42: -0.46307635
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbf874a2f; // action43: -1.05695140
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3ec9c3a3; // action44:  0.39407071
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3f8b11ea; // action45:  1.08648419
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h3f66bdd6; // action46:  0.90133417
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3b81a4b0; // action47:  0.00395640
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'hbfb95963; // action48: -1.44804037
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbfce31a2; // action49: -1.61088967
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h3f87942f; // action50:  1.05920970
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbfd90549; // action51: -1.69547379
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbfcf406c; // action52: -1.61915350
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h3fa95ed4; // action53:  1.32320642
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3f0541bf; // action54:  0.52053446
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h3f81fb6a; // action55:  1.01548505
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'hbfbf2bff; // action56: -1.49353015
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbe486840; // action57: -0.19571018
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'hbf1cc01d; // action58: -0.61230642
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'hbdefdc79; // action59: -0.11711974
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbedf1240; // action60: -0.43568611
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'hbf3c7154; // action61: -0.73610425
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'hbff352b2; // action62: -1.90096116
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3fd6eba4; // action63:  1.67906618
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3eea80d4; // action64:  0.45801413
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'hbf57d23d; // action65: -0.84305173
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h3fd8b62c; // action66:  1.69305944
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h3f917124; // action67:  1.13626528
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'hbfbd9b8a; // action68: -1.48130918
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'hbe9fb94e; // action69: -0.31196064
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h3ffc881d; // action70:  1.97290385
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3f98fcb7; // action71:  1.19521224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'hbe473acd; // action72: -0.19456024
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3fac8216; // action73:  1.34771991
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'hbf37d0c8; // action74: -0.71802950
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3f87e3c1; // action75:  1.06163800
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h3e05051c; // action76:  0.12990230
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h3eef3ff6; // action77:  0.46728486
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbfd403fb; // action78: -1.65637147
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbea8447a; // action79: -0.32864743
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3faa1092; // action80:  1.32863069
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3fd3a7d3; // action81:  1.65355909
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h3fa20802; // action82:  1.26586938
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'hbebd6157; // action83: -0.36988327
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbf253e50; // action84: -0.64548206
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbfb9733b; // action85: -1.44882905
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h3fdcc720; // action86:  1.72482681
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3fb872c5; // action87:  1.44100249
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbe108300; // action88: -0.14112473
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h3e62431b; // action89:  0.22095911
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'hbdad5624; // action90: -0.08463696
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'hbe22b4b8; // action91: -0.15889251
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h3f443b48; // action92:  0.76652956
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h3f458adb; // action93:  0.77165002
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'hbf0a3024; // action94: -0.53979707
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h3f84e5cc; // action95:  1.03826284
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h3f71545e; // action96:  0.94269359
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3b4232c0; // action97:  0.00296323
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h3fbd7b3f; // action98:  1.48032367
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3f87023d; // action99:  1.05475581
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'hbfacbae4; // action100: -1.34945345
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'hbf960f07; // action101: -1.17233360
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3f916c8f; // action102:  1.13612545
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbffa2292; // action103: -1.95418000
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h3fe11a1d; // action104:  1.75860941
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbf73603e; // action105: -0.95068729
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'hbf9e942a; // action106: -1.23889661
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h3f5ec6a3; // action107:  0.87021846
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'hbf9856a1; // action108: -1.19014370
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3fa78dd4; // action109:  1.30901575
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h3fbb6ae3; // action110:  1.46419942
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbf989c88; // action111: -1.19227695
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3e138eb3; // action112:  0.14409904
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'hbf6a33dc; // action113: -0.91485381
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'hbe8585cd; // action114: -0.26078644
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'hbff19644; // action115: -1.88739824
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'hbcfe6d33; // action116: -0.03105793
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'hbf777b78; // action117: -0.96672773
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3f73b389; // action118:  0.95195824
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3fd1df79; // action119:  1.63963234
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'hbfbfe0ad; // action120: -1.49904406
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'hbfe946e0; // action121: -1.82247543
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'hbf8a4e80; // action122: -1.08052063
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3f4888d3; // action123:  0.78333777
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'hbf0e581d; // action124: -0.55603200
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h3fa1da0c; // action125:  1.26446676
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbf3166d5; // action126: -0.69297534
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3fbec68d; // action127:  1.49043429
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h3f7c34b1; // action128:  0.98517901
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3ed34cde; // action129:  0.41269583
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'hbf887c3b; // action130: -1.06629121
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h3fe8803f; // action131:  1.81641376
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'hbfdac78e; // action132: -1.70921493
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'hbecd74a7; // action133: -0.40128061
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'hbffa8b1d; // action134: -1.95737040
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h3f0d3d58; // action135:  0.55171728
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'hbfaf7a62; // action136: -1.37092233
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'hbf1a8ca7; // action137: -0.60370868
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h3fa844bc; // action138:  1.31459761
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h3f083122; // action139:  0.53199971
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'hbfa74426; // action140: -1.30676723
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h3fe02bad; // action141:  1.75133288
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3f9fff51; // action142:  1.24997914
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'hbf946848; // action143: -1.15943241
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'hbf5f97f0; // action144: -0.87341213
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h3f768634; // action145:  0.96298528
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'hbf67d408; // action146: -0.90557909
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbf6f3bfa; // action147: -0.93450892
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'hbfd65c8b; // action148: -1.67469919
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbf963fb1; // action149: -1.17381871
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h3f10d985; // action150:  0.56581908
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h3f51189d; // action151:  0.81678182
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'hbf9b6312; // action152: -1.21396089
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3fef8869; // action153:  1.87135041
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'hbf1fce64; // action154: -0.62424302
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h3ed93a6d; // action155:  0.42427388
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbe652efb; // action156: -0.22381203
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h3feb028b; // action157:  1.83601511
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbec3b281; // action158: -0.38222125
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'hbf62bd20; // action159: -0.88569832
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbfbdfcc5; // action160: -1.48427641
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'hbf2373c7; // action161: -0.63848537
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h3f81a69a; // action162:  1.01289678
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h3f3b8bdc; // action163:  0.73260283
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbec43a78; // action164: -0.38325858
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3f412c90; // action165:  0.75458622
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbfd51e3a; // action166: -1.66498494
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h3ed9cfaf; // action167:  0.42541263
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3f663274; // action168:  0.89920735
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbeaefcce; // action169: -0.34177250
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbe13628a; // action170: -0.14393058
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3fb78015; // action171:  1.43359625
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'hbfb17c6a; // action172: -1.38660932
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3ed4f7ab; // action173:  0.41595206
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'hbf26b060; // action174: -0.65112877
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3f02e5eb; // action175:  0.51132077
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3fa81d52; // action176:  1.31339478
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h3fd21655; // action177:  1.64130652
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbf56708e; // action178: -0.83765495
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h3fc0779f; // action179:  1.50365055
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h3f7fe7ee; // action180:  0.99963272
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbd5fef26; // action181: -0.05467143
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h3f894ffc; // action182:  1.07275343
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h3e8cbe47; // action183:  0.27488920
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'hbfb0d76d; // action184: -1.38157427
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h3ffeffef; // action185:  1.99218547
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3fdd533b; // action186:  1.72910249
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'hbfb03d35; // action187: -1.37686789
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbf63049c; // action188: -0.88678908
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbf5079d4; // action189: -0.81435895
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'hbf91af24; // action190: -1.13815737
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'hbe2b4cf4; // action191: -0.16728574

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 11:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbfe755f2; // action0: -1.80731034
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'hbfa193d4; // action1: -1.26232386
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3f9d995e; // action2:  1.23124290
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'hbfa118b8; // action3: -1.25856686
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3db5d4da; // action4:  0.08878489
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbe59050f; // action5: -0.21193336
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3fca8284; // action6:  1.58210802
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbffad43b; // action7: -1.95960176
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'hbfa3353d; // action8: -1.27506220
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbf9e47ca; // action9: -1.23656583
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'hbf49546e; // action10: -0.78644454
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbf585100; // action11: -0.84498596
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'hbf2e2824; // action12: -0.68030000
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbfc649da; // action13: -1.54912877
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbf21b530; // action14: -0.63167095
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3fbee5fd; // action15:  1.49139369
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h3f6d82d0; // action16:  0.92777729
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'hbfa5aa5a; // action17: -1.29426122
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'hbf70ce63; // action18: -0.94064921
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbf089345; // action19: -0.53349715
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h3c100a44; // action20:  0.00879151
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h3ecb4b53; // action21:  0.39705905
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'hbf10ee8c; // action22: -0.56613994
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbfd4342b; // action23: -1.65784204
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h3fdee689; // action24:  1.74141037
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'hbfca3ba1; // action25: -1.57994473
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h3fef555a; // action26:  1.86979222
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'hbed64854; // action27: -0.41852057
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'hbfafe9ab; // action28: -1.37431848
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h3f9abd3c; // action29:  1.20889997
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'hbfd6c503; // action30: -1.67788732
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbfcc15bd; // action31: -1.59441340
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbf78cf3c; // action32: -0.97191215
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'hbe2d9dcc; // action33: -0.16954726
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'hbe870bc7; // action34: -0.26376173
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3f087783; // action35:  0.53307360
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'hbfef8e9e; // action36: -1.87153983
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h3e946d06; // action37:  0.28989428
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbfed8183; // action38: -1.85551488
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'hbea98a93; // action39: -0.33113536
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3ff26e4d; // action40:  1.89399111
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbdbdd76d; // action41: -0.09269605
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3fa28a9d; // action42:  1.26985514
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h3f025e90; // action43:  0.50925541
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'hbde38d66; // action44: -0.11110954
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3e545af6; // action45:  0.20737824
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h3ff26d8f; // action46:  1.89396846
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3fea8ae6; // action47:  1.83236384
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h3fb53ac3; // action48:  1.41585577
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h3f890208; // action49:  1.07037449
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h3f37aacb; // action50:  0.71744984
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbe2706a8; // action51: -0.16311133
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h3f7d0e81; // action52:  0.98850256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'hbfb11de5; // action53: -1.38372481
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3fa5c381; // action54:  1.29502881
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'hbf56fe1b; // action55: -0.83981484
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'hbfc4f28f; // action56: -1.53865230
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h3f29fb0b; // action57:  0.66398686
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3fca4405; // action58:  1.58020079
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h3eb9c756; // action59:  0.36284894
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbf2b3d70; // action60: -0.66890621
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'hbf87b7ff; // action61: -1.06030262
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'hbfdf14fc; // action62: -1.74282789
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'hbf832f1a; // action63: -1.02487493
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3fa88925; // action64:  1.31668532
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3ee47487; // action65:  0.44620153
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbe4cac1d; // action66: -0.19987531
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbd823c5f; // action67: -0.06359171
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'hbebfdd6f; // action68: -0.37473628
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3fe8e47e; // action69:  1.81947303
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'hbe8ac304; // action70: -0.27101910
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'hbfa6b14d; // action71: -1.30228579
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3f0bbe9a; // action72:  0.54587710
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3f4a1a31; // action73:  0.78946215
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'hbf61424a; // action74: -0.87991774
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3f876a6d; // action75:  1.05793536
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'hbf8f35ac; // action76: -1.11882544
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h3e41b2c3; // action77:  0.18915848
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbff8f7ef; // action78: -1.94506633
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h3cd4f1d5; // action79:  0.02599422
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3fb1b475; // action80:  1.38831961
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'hbfe4477b; // action81: -1.78343141
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h3efab9f7; // action82:  0.48970005
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'hbf59a9ee; // action83: -0.85024917
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h3e79fa31; // action84:  0.24411847
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbf83f1c8; // action85: -1.03081608
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'hbf86fea8; // action86: -1.05464649
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3f99f83c; // action87:  1.20288801
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h3fe363b5; // action88:  1.77648032
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbfb1daf0; // action89: -1.38949394
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3f0ff702; // action90:  0.56236279
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'hbf69f429; // action91: -0.91388184
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbe4621c4; // action92: -0.19348818
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'hbfd634d0; // action93: -1.67348671
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3f10388e; // action94:  0.56336296
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h3fa6e42b; // action95:  1.30383813
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'hbe0a00c8; // action96: -0.13476861
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3f87b65e; // action97:  1.06025290
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbfedc5ba; // action98: -1.85759664
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'hbfdc6510; // action99: -1.72183418
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h3fadcfdc; // action100:  1.35790586
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'hbeed1fff; // action101: -0.46313474
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3f96b65d; // action102:  1.17744029
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbf6bcf42; // action103: -0.92113125
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'hbeb277ac; // action104: -0.34856927
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbf979f46; // action105: -1.18454814
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3f545dde; // action106:  0.82955730
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h3e16f68e; // action107:  0.14742491
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3fae4398; // action108:  1.36143780
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3ed484c5; // action109:  0.41507545
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'hbedf443e; // action110: -0.43606752
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h3fd9ae41; // action111:  1.70063031
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3fe6339d; // action112:  1.79845011
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'hbfdb9f59; // action113: -1.71580040
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h3fc62aa1; // action114:  1.54817593
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3fa14b2f; // action115:  1.26010692
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'hbf8d2946; // action116: -1.10282207
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3ddec633; // action117:  0.10877647
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'hbf39d0d7; // action118: -0.72584289
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3f51402b; // action119:  0.81738538
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h3f146c03; // action120:  0.57977313
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'hbeef36ce; // action121: -0.46721500
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'hbf258fe0; // action122: -0.64672661
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3faaa508; // action123:  1.33316135
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'hbf44ac93; // action124: -0.76825827
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h3f68184f; // action125:  0.90662092
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbe59fc27; // action126: -0.21287595
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3ec2fc09; // action127:  0.38082913
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'hbf13af43; // action128: -0.57689303
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3f64437f; // action129:  0.89165491
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'hbe06d4f1; // action130: -0.13167168
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbf81abc6; // action131: -1.01305461
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'hbec52f23; // action132: -0.38512525
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'hbe92d334; // action133: -0.28676760
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'hbf99bbc8; // action134: -1.20104313
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h3e3b8e26; // action135:  0.18315944
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'hbfbbf1b1; // action136: -1.46831334
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h3e03434a; // action137:  0.12818637
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'hbfd4270b; // action138: -1.65744150
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'hbfee15a5; // action139: -1.86003554
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h3fce7aad; // action140:  1.61311877
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'hbfc2657d; // action141: -1.51872218
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'hbe6a8102; // action142: -0.22900775
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'hbf925221; // action143: -1.14313138
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'hbf4fcd97; // action144: -0.81173080
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'hbdcaba76; // action145: -0.09898846
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h3fd64f10; // action146:  1.67428780
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h3fd4bd89; // action147:  1.66203415
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'hbf281093; // action148: -0.65650290
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h3fec3fe4; // action149:  1.84569979
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h3ed48a3b; // action150:  0.41511711
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h3fa2f081; // action151:  1.27296460
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3fd2fc90; // action152:  1.64833260
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'hbfe005df; // action153: -1.75017917
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'hbe02491f; // action154: -0.12723206
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'hbfa6011e; // action155: -1.29690909
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbe6d5f74; // action156: -0.23180944
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h3ed81c71; // action157:  0.42209199
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h3f20171b; // action158:  0.62535256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h3fe2fea4; // action159:  1.77339602
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h3fc43b21; // action160:  1.53305447
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'hbff1308f; // action161: -1.88429439
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h3eae626c; // action162:  0.34059465
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h3f8e6dc0; // action163:  1.11272430
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h3fcffe31; // action164:  1.62494481
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3fc06ebf; // action165:  1.50337970
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h3f9d3780; // action166:  1.22825623
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbeb58dbc; // action167: -0.35459697
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'hbff12871; // action168: -1.88404667
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbfddf1c7; // action169: -1.73394096
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h3fec9b04; // action170:  1.84848070
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3f8eede9; // action171:  1.11663544
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3f548327; // action172:  0.83012623
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3f3e7855; // action173:  0.74402362
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3db599a8; // action174:  0.08867198
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'hbdd30a2d; // action175: -0.10304675
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3eece61b; // action176:  0.46269307
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'hbf26fbcd; // action177: -0.65227968
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbfa298ac; // action178: -1.27028418
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbfc08d33; // action179: -1.50430906
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'hbd8b89c0; // action180: -0.06813383
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbf8a0db8; // action181: -1.07854366
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbf579313; // action182: -0.84208792
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h3eda80b2; // action183:  0.42676312
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3fadc2ac; // action184:  1.35750341
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbd91f3b8; // action185: -0.07126564
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3e3a3255; // action186:  0.18183263
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h3ff41145; // action187:  1.90677702
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbfcd3934; // action188: -1.60330820
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h3e9c68cc; // action189:  0.30548704
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'hbf4e45d0; // action190: -0.80575275
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h3f207e5c; // action191:  0.62692809

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 12:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbfc0bbfb; // action0: -1.50573671
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3fe83fe4; // action1:  1.81444979
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'hbf5ec8d9; // action2: -0.87025219
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3ff7cf6d; // action3:  1.93601763
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3fa9054d; // action4:  1.32047427
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbfa5f875; // action5: -1.29664481
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'hbfb9eea0; // action6: -1.45259476
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbf92cb25; // action7: -1.14682448
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'hbee2d2cc; // action8: -0.44301450
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbf9d76ff; // action9: -1.23019397
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h3fc18fe5; // action10:  1.51220381
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h3d454636; // action11:  0.04816266
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h3f048dda; // action12:  0.51778948
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbee7fbf2; // action13: -0.45309407
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbfa4912c; // action14: -1.28568029
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3fcd09ee; // action15:  1.60186553
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h3fbc5c44; // action16:  1.47156572
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h3fe6a3a6; // action17:  1.80186915
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'hbeed66b4; // action18: -0.46367419
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h3f3710a0; // action19:  0.71509743
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'hbf4068bb; // action20: -0.75159806
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbe884a83; // action21: -0.26619348
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'hbf44f083; // action22: -0.76929492
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbfbcd7fd; // action23: -1.47534144
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbe0e71cb; // action24: -0.13910596
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'hbfc098e8; // action25: -1.50466633
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'hbfb72775; // action26: -1.43089163
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'hbf10614a; // action27: -0.56398451
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3fdfe7d4; // action28:  1.74926233
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h3f98a1bf; // action29:  1.19243610
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'hbfecf8c5; // action30: -1.85134184
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbf9148c9; // action31: -1.13503373
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbda0f117; // action32: -0.07858484
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3fdde79e; // action33:  1.73363090
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h3f71d0cc; // action34:  0.94459224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'hbfaefc33; // action35: -1.36707151
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'hbfe7c4c0; // action36: -1.81069183
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'hbf81fc0a; // action37: -1.01550412
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h3fffef79; // action38:  1.99949563
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'hbfdae5f5; // action39: -1.71014273
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3f81eec8; // action40:  1.01509953
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbe525349; // action41: -0.20539583
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3ed22a49; // action42:  0.41047886
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbee53e90; // action43: -0.44774294
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3dfc6d83; // action44:  0.12325575
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3f9b40da; // action45:  1.21291661
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbb9bc808; // action46: -0.00475407
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'hbfb34db4; // action47: -1.40080881
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'hbf8dfed5; // action48: -1.10933936
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h3e9732b1; // action49:  0.29530862
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbf88e370; // action50: -1.06944084
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbf8c1da3; // action51: -1.09465444
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbf9020d4; // action52: -1.12600183
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h3fe5c129; // action53:  1.79495728
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'hbf9663dd; // action54: -1.17492259
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'hbff47a2f; // action55: -1.90997875
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'hbf4f51f6; // action56: -0.80984437
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbfce6c7c; // action57: -1.61268568
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'hbfbdb40a; // action58: -1.48205686
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h3f3be641; // action59:  0.73398215
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbf4782d4; // action60: -0.77934003
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3d696e43; // action61:  0.05698992
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3f0b8142; // action62:  0.54494107
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'hbe18adc7; // action63: -0.14910041
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'hbf5e6263; // action64: -0.86868876
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3fee6e83; // action65:  1.86274755
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbfaf179c; // action66: -1.36790800
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h3ec580a4; // action67:  0.38574708
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3e40c33c; // action68:  0.18824476
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'hbf74e7c4; // action69: -0.95666146
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'hbf46a01a; // action70: -0.77588046
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'hbf5a4e37; // action71: -0.85275596
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3ef7737c; // action72:  0.48330295
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3f6d283b; // action73:  0.92639512
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3f3a612c; // action74:  0.72804523
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3e53920b; // action75:  0.20661180
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'hbe1167a0; // action76: -0.14199686
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h3dfe73ad; // action77:  0.12424407
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h3e6cd4cb; // action78:  0.23128049
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbf89f4d2; // action79: -1.07778382
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3f3753ee; // action80:  0.71612442
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'hbe3e2e9a; // action81: -0.18572465
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h3e2af117; // action82:  0.16693531
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h3f267452; // action83:  0.65021241
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbf192e6d; // action84: -0.59836465
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbffd766a; // action85: -1.98017621
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h3e84a8e6; // action86:  0.25910109
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'hbfa3f492; // action87: -1.28090119
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbfa4ee4f; // action88: -1.28852260
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h3ffec867; // action89:  1.99049079
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3eb2992c; // action90:  0.34882486
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'hbf856d09; // action91: -1.04238999
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h3fbf852c; // action92:  1.49625158
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'hbfe4bd2a; // action93: -1.78702283
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3f792bd3; // action94:  0.97332495
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h3fd5cd60; // action95:  1.67033005
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'hbed5b062; // action96: -0.41736132
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'hbeea28b7; // action97: -0.45734188
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h3f1b67aa; // action98:  0.60705054
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3fef7597; // action99:  1.87077606
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'hbf9a6539; // action100: -1.20621407
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h3de9e8ae; // action101:  0.11421333
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3e0164cd; // action102:  0.12636109
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h3fb602cc; // action103:  1.42196035
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h3f95a686; // action104:  1.16914439
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbfdabcc9; // action105: -1.70888627
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'hbe2bff97; // action106: -0.16796719
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbf9f991a; // action107: -1.24685979
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'hbfac5476; // action108: -1.34632754
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'hbecf5f45; // action109: -0.40502372
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'hbf2f5a09; // action110: -0.68496758
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbef313a2; // action111: -0.47475916
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3f51791e; // action112:  0.81825435
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'hbff2938d; // action113: -1.89512789
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h3f070437; // action114:  0.52740806
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3f8ea632; // action115:  1.11444688
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3fbfd629; // action116:  1.49872315
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3f5d024e; // action117:  0.86331642
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3f3e922e; // action118:  0.74441803
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3fecda4a; // action119:  1.85041165
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'hbff86dc6; // action120: -1.94085002
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'hbffd876e; // action121: -1.98069549
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'hbf5e92fe; // action122: -0.86943042
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'hbfd3e15c; // action123: -1.65531492
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3f1c5740; // action124:  0.61070633
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'hbead1e95; // action125: -0.33812395
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h3fafb624; // action126:  1.37274599
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3faf79d9; // action127:  1.37090600
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'hbf92f921; // action128: -1.14822781
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'hbf6d909c; // action129: -0.92798781
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h3f649903; // action130:  0.89295977
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h3ffbc23b; // action131:  1.96686494
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h3fd9b5c8; // action132:  1.70086002
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'hbf977a8b; // action133: -1.18342721
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3ffd88f1; // action134:  1.98074162
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'hbd8c6e7c; // action135: -0.06857011
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h3f270b2a; // action136:  0.65251410
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'hbf8a5a4e; // action137: -1.08088088
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'hbfe12557; // action138: -1.75895202
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h3e5ae0d5; // action139:  0.21374829
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h3f0939ff; // action140:  0.53604120
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'hbf373357; // action141: -0.71562713
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3e5d2565; // action142:  0.21596296
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'hbfaf807b; // action143: -1.37110841
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'hbe285810; // action144: -0.16439843
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'hbfa33845; // action145: -1.27515471
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'hbeeb6807; // action146: -0.45977804
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbf9df45d; // action147: -1.23401988
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3f357f67; // action148:  0.70897526
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h3f9ec6b9; // action149:  1.24043953
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h3fd608bb; // action150:  1.67214143
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbe8fba01; // action151: -0.28071597
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3dbcbba0; // action152:  0.09215474
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3fd0f2b4; // action153:  1.63240671
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h3e1cef62; // action154:  0.15325692
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'hbeb4ec8a; // action155: -0.35336715
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbfc194c3; // action156: -1.51235235
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h3fde2abd; // action157:  1.73567927
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbf5d6349; // action158: -0.86479622
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'hbfb326fd; // action159: -1.39962733
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbf9b20c5; // action160: -1.21193755
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'hbeef6371; // action161: -0.46755555
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'hbf8c459f; // action162: -1.09587467
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'hbf7ff8d7; // action163: -0.99989074
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbfa81308; // action164: -1.31308079
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3fabecd6; // action165:  1.34316516
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbe9ed957; // action166: -0.31025192
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h3fb72dd2; // action167:  1.43108582
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'hbede5791; // action168: -0.43426183
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h3f8eb62f; // action169:  1.11493480
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h3fd52333; // action170:  1.66513669
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'hbf0da361; // action171: -0.55327421
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3fd50735; // action172:  1.66428244
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'hbfb6d654; // action173: -1.42841578
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'hbf8f4e9a; // action174: -1.11958623
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3f5e1276; // action175:  0.86746919
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3fd001d4; // action176:  1.62505579
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h3d402f0d; // action177:  0.04691987
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbfdc1f3e; // action178: -1.71970344
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h3ed40b17; // action179:  0.41414711
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h3f960939; // action180:  1.17215645
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbf0a85be; // action181: -0.54110324
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h3eb3ebe1; // action182:  0.35140899
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'hbefce756; // action183: -0.49395245
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3f021471; // action184:  0.50812441
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbf2b44a6; // action185: -0.66901624
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'hbfbcd681; // action186: -1.47529614
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h3d9217d3; // action187:  0.07133450
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbeb5b635; // action188: -0.35490575
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h3f565cce; // action189:  0.83735359
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'hbf184de5; // action190: -0.59493858
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'hbfca97f2; // action191: -1.58276200

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 13:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbfb093df; // action0: -1.37951267
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'hbfbb8c61; // action1: -1.46522152
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3e8e8023; // action2:  0.27832136
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3f88308f; // action3:  1.06398189
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3fb84b75; // action4:  1.43980277
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h3f9829c6; // action5:  1.18877482
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'hbf80c459; // action6: -1.00599205
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h3be907ab; // action7:  0.00711151
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'hbd1c9ed7; // action8: -0.03823742
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbf5aa72b; // action9: -0.85411328
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'hbe9f0c4b; // action10: -0.31064066
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h3eefe000; // action11:  0.46850586
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h3f0bf5ec; // action12:  0.54672122
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbff764e4; // action13: -1.93276644
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbfbc3ac7; // action14: -1.47054374
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3e62fea8; // action15:  0.22167456
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'hbf592fab; // action16: -0.84838361
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'hbf86d41e; // action17: -1.05334830
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'hbfd98c7e; // action18: -1.69959998
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbee56ce1; // action19: -0.44809631
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'hbfeb0668; // action20: -1.83613300
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbfda295a; // action21: -1.70438695
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h3fb25cca; // action22:  1.39345670
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h3f7c453b; // action23:  0.98543137
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'h3e837799; // action24:  0.25677183
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'hbfe9ada2; // action25: -1.82561135
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h3f10e730; // action26:  0.56602764
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'hbf8eeba2; // action27: -1.11656594
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'hbf06098b; // action28: -0.52358311
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbf78b037; // action29: -0.97143883
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'hbfd1b33e; // action30: -1.63828254
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbfa9864a; // action31: -1.32441068
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbf1fc336; // action32: -0.62407243
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3fb2fbcb; // action33:  1.39830911
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'hbfa13a52; // action34: -1.25959229
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3ebec719; // action35:  0.37261274
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3d535420; // action36:  0.05159390
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'hbfdc03b3; // action37: -1.71886289
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h3f499461; // action38:  0.78742033
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'hbd43f365; // action39: -0.04783954
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'hbff41215; // action40: -1.90680182
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h3f221e1a; // action41:  0.63327181
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'hbf5569ee; // action42: -0.83364761
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h3fecc305; // action43:  1.84970152
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'hbfacc225; // action44: -1.34967482
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'hbfec2dfc; // action45: -1.84515333
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbf8b0af2; // action46: -1.08627152
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'hbff1f8d5; // action47: -1.89040625
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h3fcd62ad; // action48:  1.60457385
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbed95217; // action49: -0.42445442
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'h3fa96db7; // action50:  1.32366073
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h3ebea8fe; // action51:  0.37238306
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h3f8a3af3; // action52:  1.07992399
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h3f2ed9a2; // action53:  0.68300831
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3fa2f8e7; // action54:  1.27322090
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'hbfee5b4d; // action55: -1.86216128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'hbf3d3bf9; // action56: -0.73919636
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'h3e865f58; // action57:  0.26244617
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3e0c8a33; // action58:  0.13724594
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h3fea6942; // action59:  1.83133721
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h3eb6b3f4; // action60:  0.35684168
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'hbf1aa51d; // action61: -0.60408193
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3f51e4da; // action62:  0.81989825
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3f95ed6c; // action63:  1.17130804
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3f398bdb; // action64:  0.72479028
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'hbfc42441; // action65: -1.53235638
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbfe6324c; // action66: -1.79840994
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbff4c348; // action67: -1.91220951
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3eb7a6f7; // action68:  0.35869572
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3f6bd5d5; // action69:  0.92123157
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'hbf5ed129; // action70: -0.87037903
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3f812fbb; // action71:  1.00926912
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3fcc2c8e; // action72:  1.59510970
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3edba196; // action73:  0.42896718
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3fbc66af; // action74:  1.47188365
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3fb91ffc; // action75:  1.44628859
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h3ff524d2; // action76:  1.91518617
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h3fc6b309; // action77:  1.55233872
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbfb50a49; // action78: -1.41437638
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h3f8491aa; // action79:  1.03569531
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3ea832f5; // action80:  0.32851377
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3f633daf; // action81:  0.88765997
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h3fb49df2; // action82:  1.41107011
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'hbfb6d0e8; // action83: -1.42825031
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbe7763ac; // action84: -0.24159116
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h3f41ec71; // action85:  0.75751406
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h3ffd16dc; // action86:  1.97726011
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3fad1077; // action87:  1.35206497
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h3e35b351; // action88:  0.17744185
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h3f435e1f; // action89:  0.76315492
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'hbf3233b2; // action90: -0.69610131
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3f2094bc; // action91:  0.62726951
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbe2cf4f4; // action92: -0.16890317
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h3f77117f; // action93:  0.96511072
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3e9b6707; // action94:  0.30352041
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h3f278c83; // action95:  0.65448779
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h3fe7cbc6; // action96:  1.81090617
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3f916b2d; // action97:  1.13608325
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h3ef55ed1; // action98:  0.47923902
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'hbf95d8ed; // action99: -1.17068255
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'hbffb4428; // action100: -1.96301746
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'hbf5cda4b; // action101: -0.86270589
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'hbf5c23ce; // action102: -0.85992134
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbfa5d548; // action103: -1.29557133
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h3fcbe34c; // action104:  1.59287405
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h3f1c3ebc; // action105:  0.61033225
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'hbf1f0e7d; // action106: -0.62131482
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h3ff33d3a; // action107:  1.90030599
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'hbfe6fbfc; // action108: -1.80456495
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3f71dff1; // action109:  0.94482332
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'hbff90627; // action110: -1.94550025
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbf188da5; // action111: -0.59591132
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3feab7b3; // action112:  1.83373106
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'hbe9008a3; // action113: -0.28131589
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'hbf33b869; // action114: -0.70203263
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3e3aca74; // action115:  0.18241292
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3e8c4c87; // action116:  0.27402136
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'hbf8a9081; // action117: -1.08253491
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'hbf428e7e; // action118: -0.75998676
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3eb4da53; // action119:  0.35322818
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h3fe6556e; // action120:  1.79948211
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3fcbe35b; // action121:  1.59287584
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'hbf63a4c0; // action122: -0.88923264
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3fcf3877; // action123:  1.61891067
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3fedf298; // action124:  1.85896587
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'hbf8ee5e6; // action125: -1.11639094
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h3d5b20b8; // action126:  0.05349800
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3f95d22d; // action127:  1.17047656
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'hbfc30ad5; // action128: -1.52376807
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3f0576c7; // action129:  0.52134365
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'hbfbcec83; // action130: -1.47596776
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbfb7e02e; // action131: -1.43652892
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h3e252905; // action132:  0.16128929
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3f6df452; // action133:  0.92950928
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3f49cd3a; // action134:  0.78828776
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'hbff24259; // action135: -1.89264977
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h3fc1d484; // action136:  1.51429796
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'hbf8b330e; // action137: -1.08749557
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'hbe874458; // action138: -0.26419330
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h3f901151; // action139:  1.12552845
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h3fea6b27; // action140:  1.83139503
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h3ff7fea8; // action141:  1.93745899
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3fd95f48; // action142:  1.69822025
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h3ed6695c; // action143:  0.41877258
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3fc46b22; // action144:  1.53451943
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'hbef0912c; // action145: -0.46985757
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'hbfb4c15f; // action146: -1.41215122
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbf68d2ae; // action147: -0.90946472
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3f5c1e14; // action148:  0.85983396
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h3faa131a; // action149:  1.32870793
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'hbfde9bd2; // action150: -1.73913026
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbff5f13a; // action151: -1.92142415
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3fec0dc2; // action152:  1.84416986
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3eb9134c; // action153:  0.36147535
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h3f9ad9a5; // action154:  1.20976698
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h3e3a1dab; // action155:  0.18175380
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbf253708; // action156: -0.64537096
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbffee980; // action157: -1.99150085
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbfe6310d; // action158: -1.79837191
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'hbde25c57; // action159: -0.11052769
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h3f522118; // action160:  0.82081747
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h3dec6bdf; // action161:  0.11544012
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'hbfbf4a81; // action162: -1.49446118
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h3feff60a; // action163:  1.87469602
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbf6a1bc4; // action164: -0.91448617
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3fa9cefb; // action165:  1.32662904
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbea761f4; // action166: -0.32691920
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbff45c18; // action167: -1.90906048
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3fb331f3; // action168:  1.39996183
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbfedc10d; // action169: -1.85745394
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h3f92c356; // action170:  1.14658618
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'hbf6e16e5; // action171: -0.93003684
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3ebc29e9; // action172:  0.36750725
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3faa2940; // action173:  1.32938385
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3ff81482; // action174:  1.93812585
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3fd459c7; // action175:  1.65898979
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'hbf1f4ae4; // action176: -0.62223649
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h3e8a89f2; // action177:  0.27058369
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbfebf5e4; // action178: -1.84344149
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbfbb1d82; // action179: -1.46183801
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'hbf9e7877; // action180: -1.23805130
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbfedbe3b; // action181: -1.85736787
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h3fbb0258; // action182:  1.46100903
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h3ea2b94c; // action183:  0.31781995
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'hbf6411c8; // action184: -0.89089632
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbf3b2901; // action185: -0.73109442
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3f654a16; // action186:  0.89566171
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h3f584696; // action187:  0.84482706
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbfe1794f; // action188: -1.76151454
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbfa42d0a; // action189: -1.28262448
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h3f684289; // action190:  0.90726525
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h3fdfe0cc; // action191:  1.74904776

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 14:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h3f6936dc; // action0:  0.91099334
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3e12a66f; // action1:  0.14321302
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'hbfc512db; // action2: -1.53963792
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'hbfc1caa5; // action3: -1.51399672
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3fa41159; // action4:  1.28177941
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h3fadf601; // action5:  1.35906994
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'hbcbaf7d3; // action6: -0.02282325
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbfdd0281; // action7: -1.72663891
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h3f8a99ed; // action8:  1.08282244
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h3f4ef3f8; // action9:  0.80841017
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'hbf5e0ccc; // action10: -0.86738276
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h3fd2be6d; // action11:  1.64643633
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'hbea45836; // action12: -0.32098550
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h3f219caf; // action13:  0.63129705
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbfdea9ec; // action14: -1.73956060
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'hbf0ba4eb; // action15: -0.54548520
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h3f905e60; // action16:  1.12788010
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h3f088d2c; // action17:  0.53340411
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h3fb34de6; // action18:  1.40081477
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbd8dd057; // action19: -0.06924503
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'hbf006ec0; // action20: -0.50168991
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbf3a2b88; // action21: -0.72722673
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h3dba50d5; // action22:  0.09097449
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h3f9c2fcf; // action23:  1.22020900
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbe3eb6db; // action24: -0.18624441
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'hbf9d3c9c; // action25: -1.22841215
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'hbf9c2b7d; // action26: -1.22007716
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3f7a8197; // action27:  0.97853988
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3f91333e; // action28:  1.13437629
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'h3fd68cd5; // action29:  1.67617285
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3eb17fb3; // action30:  0.34667739
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbf96c25d; // action31: -1.17780650
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbd717b55; // action32: -0.05895551
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3eb7d4e2; // action33:  0.35904604
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h3edf5268; // action34:  0.43617558
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3fd4752c; // action35:  1.65982580
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3f3267e1; // action36:  0.69689757
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h3e8beba4; // action37:  0.27328217
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbfde4cc6; // action38: -1.73671794
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h3f9636dd; // action39:  1.17354929
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'hbed65623; // action40: -0.41862592
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbf823a94; // action41: -1.01741266
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'hbe7fb41e; // action42: -0.24971053
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbe545927; // action43: -0.20737134
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3faa9872; // action44:  1.33277726
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3f720206; // action45:  0.94534338
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbfab2798; // action46: -1.33714581
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3faaf355; // action47:  1.33555090
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'hbe8d8b0b; // action48: -0.27645144
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h3f500b4f; // action49:  0.81267256
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbfb7f405; // action50: -1.43713439
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbf2d6831; // action51: -0.67737108
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h3f802146; // action52:  1.00101542
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'hbe820727; // action53: -0.25396082
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3f98c455; // action54:  1.19349158
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h3fe7e0cb; // action55:  1.81154764
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h3f3328e5; // action56:  0.69984275
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbedc1ae1; // action57: -0.42989257
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3fb133cd; // action58:  1.38439333
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h3ffeb7a1; // action59:  1.98997891
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbfe0ab1f; // action60: -1.75522220
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3f9f56fd; // action61:  1.24484217
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3ffd58f7; // action62:  1.97927749
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3ffa9ea4; // action63:  1.95796633
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'hbd2018ed; // action64: -0.03908627
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'hbff1a20c; // action65: -1.88775778
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbfb6a2c8; // action66: -1.42684269
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbfe8f192; // action67: -1.81987214
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3f3172f6; // action68:  0.69316041
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3fc3acf0; // action69:  1.52871513
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h3f3e1a35; // action70:  0.74258739
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3feaf2b9; // action71:  1.83553231
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3f253f3e; // action72:  0.64549625
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3f7616b0; // action73:  0.96128368
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3f36b2a5; // action74:  0.71366340
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'hbd4a72ad; // action75: -0.04942577
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'hbf210083; // action76: -0.62891406
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbfa6e8fe; // action77: -1.30398536
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbfec818a; // action78: -1.84770322
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbf21f121; // action79: -0.63258559
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3e3bffb7; // action80:  0.18359266
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'hbff40e09; // action81: -1.90667832
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'hbecd2a74; // action82: -0.40071452
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'hbc8c11f7; // action83: -0.01709841
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h3f0050b4; // action84:  0.50123143
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbf975425; // action85: -1.18225539
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'hbeaf3f27; // action86: -0.34227869
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'hbff1787b; // action87: -1.88648927
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'h3fe534d7; // action88:  1.79067504
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbe9debfe; // action89: -0.30844110
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'hbfbd4881; // action90: -1.47877514
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'hbe8e0494; // action91: -0.27737868
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbe274c33; // action92: -0.16337661
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h3fd6bb16; // action93:  1.67758441
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'hbf8ddfc8; // action94: -1.10839176
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'hbf46428a; // action95: -0.77445281
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h3f917a22; // action96:  1.13653970
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3f9ca9ab; // action97:  1.22392786
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbc5847aa; // action98: -0.01320068
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'hbff763b5; // action99: -1.93273032
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'hbfcb09f3; // action100: -1.58624113
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'hbea58e75; // action101: -0.32335249
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3ff082ec; // action102:  1.87899542
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h3f6d16dc; // action103:  0.92613006
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h3fe1f592; // action104:  1.76530671
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbf902c9d; // action105: -1.12636149
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'hbf6284a5; // action106: -0.88483649
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbf4469a7; // action107: -0.76723713
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3f98194a; // action108:  1.18827176
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3ff0787f; // action109:  1.87867725
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h3fa1875e; // action110:  1.26194358
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbfa81417; // action111: -1.31311309
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3f64b890; // action112:  0.89344120
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h3fa619df; // action113:  1.29766452
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'hbee170a2; // action114: -0.44031245
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3f43cc2e; // action115:  0.76483428
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'hbe591a51; // action116: -0.21201445
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3f048179; // action117:  0.51760060
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'hbfad08d1; // action118: -1.35183156
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3fcfe59c; // action119:  1.62419462
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'hbf53aa89; // action120: -0.82682091
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3fb7c841; // action121:  1.43579876
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h3fe315e2; // action122:  1.77410531
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3face17a; // action123:  1.35063100
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3f01d66b; // action124:  0.50717801
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'h3fcdf350; // action125:  1.60898781
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbf53725e; // action126: -0.82596385
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3f9dc927; // action127:  1.23270118
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'hbeafea85; // action128: -0.34358612
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'hbe6f2af5; // action129: -0.23356231
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h3f0e6a29; // action130:  0.55630738
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbef3b4ba; // action131: -0.47598821
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'hbf6f9605; // action132: -0.93588287
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'hbd8cdf3b; // action133: -0.06878515
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3fe82b57; // action134:  1.81382263
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'hbfe114c3; // action135: -1.75844610
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h3fe55a75; // action136:  1.79182303
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h3fd6cb39; // action137:  1.67807686
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h3fd77c08; // action138:  1.68347263
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h3ea74647; // action139:  0.32670805
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'hbfc8d687; // action140: -1.56904685
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'hbf577d3d; // action141: -0.84175473
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3e1bbdc4; // action142:  0.15209109
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'hbf453158; // action143: -0.77028418
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3f5a9ae4; // action144:  0.85392594
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'hbeaae8e0; // action145: -0.33380795
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h3ff37344; // action146:  1.90195513
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbe72e28d; // action147: -0.23719235
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3f9ac824; // action148:  1.20923281
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbfa9b984; // action149: -1.32597399
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'hbfc02e60; // action150: -1.50141525
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbec94606; // action151: -0.39311236
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3e8ba204; // action152:  0.27272046
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'hbfa4bda5; // action153: -1.28703749
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h3e6efcab; // action154:  0.23338573
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h3fd92f36; // action155:  1.69675326
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbf7b9751; // action156: -0.98277766
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h3e0d2254; // action157:  0.13782626
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbeb83da9; // action158: -0.35984543
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h3fcf4dfb; // action159:  1.61956728
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbf8e3f67; // action160: -1.11130989
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'hbfb0dbb5; // action161: -1.38170493
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h3f7303de; // action162:  0.94927776
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h3fdc0453; // action163:  1.71888196
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbf17fab0; // action164: -0.59366894
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3f512fbe; // action165:  0.81713474
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbd9f421a; // action166: -0.07776280
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbff3c921; // action167: -1.90457547
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3f9a1f8f; // action168:  1.20408809
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h3fd0d4b9; // action169:  1.63149178
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbf86e22b; // action170: -1.05377710
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'hbf50b9cf; // action171: -0.81533521
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3f102745; // action172:  0.56309921
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3f28813b; // action173:  0.65822190
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3f813985; // action174:  1.00956786
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'hbf0c704e; // action175: -0.54858863
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3ffd835a; // action176:  1.98057103
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'h3df169a7; // action177:  0.11787730
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbff4bbed; // action178: -1.91198504
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbea004cd; // action179: -0.31253663
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h3ff6070d; // action180:  1.92209017
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbed88d08; // action181: -0.42295098
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbe43dda6; // action182: -0.19127521
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'hbfa9be9e; // action183: -1.32612967
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3ec9d41c; // action184:  0.39419639
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'h3ff311d5; // action185:  1.89898169
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3f5bb14b; // action186:  0.85817403
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h3d44fcbf; // action187:  0.04809260
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbb94d77d; // action188: -0.00454229
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbe9e557b; // action189: -0.30924591
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h3f133ca3; // action190:  0.57514399
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'hbfcbbcfc; // action191: -1.59170485

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 15:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbd90c504; // action0: -0.07068828
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3fa9f769; // action1:  1.32786286
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3f83c161; // action2:  1.02933896
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3f9f8523; // action3:  1.24625051
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'hbecece92; // action4: -0.40391976
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h3fb03f49; // action5:  1.37693131
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3e1ee255; // action6:  0.15516026
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h3ff90c22; // action7:  1.94568276
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h3f86920b; // action8:  1.05133188
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h3f1d994f; // action9:  0.61562055
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'hbfb45710; // action10: -1.40890694
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbfdb7ab2; // action11: -1.71468186
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h3e7ab4bc; // action12:  0.24483007
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h3f427d0d; // action13:  0.75972062
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbf4ff185; // action14: -0.81227905
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'hbdd61bd5; // action15: -0.10454527
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h3fb6dbeb; // action16:  1.42858636
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'hbf7afb60; // action17: -0.98039818
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h3e386b7e; // action18:  0.18009755
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h3f6f0fa5; // action19:  0.93383247
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h3ffe302e; // action20:  1.98584533
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h3fc24ce9; // action21:  1.51797211
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h3faeb979; // action22:  1.36503518
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbdae3f62; // action23: -0.08508183
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbec778b7; // action24: -0.38959286
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'hbe8f59f3; // action25: -0.27998313
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'hbf3d4330; // action26: -0.73930645
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3f64db84; // action27:  0.89397454
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3ff136f6; // action28:  1.88448977
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbe2ddd96; // action29: -0.16979060
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'hbf8d9136; // action30: -1.10599399
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbfb62af2; // action31: -1.42318559
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbfed5a51; // action32: -1.85431874
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'hbe8e981a; // action33: -0.27850419
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h3f996026; // action34:  1.19824672
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3f965701; // action35:  1.17453015
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'hbffed9fe; // action36: -1.99102759
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h3f8272ff; // action37:  1.01913440
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbf2c35d6; // action38: -0.67269647
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'hbeee35ff; // action39: -0.46525571
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3eb8d349; // action40:  0.36098698
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbc84c3ea; // action41: -0.01620670
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3e9bc42a; // action42:  0.30423099
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbf867a16; // action43: -1.05060077
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3ed744ee; // action44:  0.42044777
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3eed0aec; // action45:  0.46297395
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h3f3f0c5a; // action46:  0.74628222
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'hbfe67d64; // action47: -1.80070162
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'hbfcd9cf9; // action48: -1.60635293
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'hbed9b3d0; // action49: -0.42519999
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbfa14247; // action50: -1.25983512
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbfe22e2d; // action51: -1.76703417
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbfec0520; // action52: -1.84390640
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h3ee4afe9; // action53:  0.44665459
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3f81dd98; // action54:  1.01457500
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'hbf8ac88d; // action55: -1.08424532
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h3fe45f9c; // action56:  1.78416777
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbfaba780; // action57: -1.34104919
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3fb51870; // action58:  1.41480827
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h3f6e8af7; // action59:  0.93180794
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h3e253850; // action60:  0.16134763
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3ffddf64; // action61:  1.98337984
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'hbeefc334; // action62: -0.46828616
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'hbf6706ca; // action63: -0.90244734
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3f1ced49; // action64:  0.61299568
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3facbc2f; // action65:  1.34949291
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbfeace07; // action66: -1.83441246
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbf74ad39; // action67: -0.95576817
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'hbfc1fcf9; // action68: -1.51553261
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'hbfa0b161; // action69: -1.25541317
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'hbf8c5800; // action70: -1.09643555
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3f020ab2; // action71:  0.50797570
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3cae6549; // action72:  0.02128853
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'hbfdb3b60; // action73: -1.71274948
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'hbf95b4a8; // action74: -1.16957569
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'hbfd56424; // action75: -1.66711855
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h3ffd2318; // action76:  1.97763348
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbf721a2f; // action77: -0.94571203
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h3eff2e85; // action78:  0.49840179
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h3f096434; // action79:  0.53668523
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3f9d6be0; // action80:  1.22985458
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3f9eb058; // action81:  1.23975658
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'h3f314be7; // action82:  0.69256443
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'hbfaa2204; // action83: -1.32916307
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h3fb96101; // action84:  1.44827282
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbf63979c; // action85: -0.88903213
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'hbc197eac; // action86: -0.00936858
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'hbfaaac61; // action87: -1.33338559
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbecbfca8; // action88: -0.39841199
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbebf7e4c; // action89: -0.37401044
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3f9187b1; // action90:  1.13695347
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'hbf185dec; // action91: -0.59518313
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbe413df3; // action92: -0.18871288
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'hbf91d5fc; // action93: -1.13934278
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'hbe95a739; // action94: -0.29229143
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'hbeed9b8a; // action95: -0.46407729
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h3eb826b1; // action96:  0.35967019
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3f347efd; // action97:  0.70506269
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbfb61fd5; // action98: -1.42284644
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'hbf908607; // action99: -1.12909019
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h3f5e71ce; // action100:  0.86892402
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h3f9c12c1; // action101:  1.21932232
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3ff05a3f; // action102:  1.87775409
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h3f1e8cbd; // action103:  0.61933500
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'hbf91ce29; // action104: -1.13910401
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h3fd5deed; // action105:  1.67086565
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3fa7e742; // action106:  1.31174493
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h3e0244d2; // action107:  0.12721565
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3f9c5d0b; // action108:  1.22158945
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3f99ec25; // action109:  1.20251906
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'hbfab26ce; // action110: -1.33712173
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbf039b96; // action111: -0.51409280
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3ff82e5f; // action112:  1.93891513
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'hbdaa749b; // action113: -0.08323022
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'hbfd9e3bc; // action114: -1.70226240
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'hbf9de333; // action115: -1.23349607
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3f436717; // action116:  0.76329178
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'hbddf467b; // action117: -0.10902115
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3f88a5ad; // action118:  1.06755602
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3f49ecfe; // action119:  0.78877246
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'hbeff2f50; // action120: -0.49840784
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'hbf9c21c5; // action121: -1.21978056
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'hbf86ba8b; // action122: -1.05256784
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3fabebc1; // action123:  1.34313214
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3f054675; // action124:  0.52060634
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'hbf870817; // action125: -1.05493438
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbf862975; // action126: -1.04814017
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'hbe84a8f9; // action127: -0.25910166
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'hbf05c855; // action128: -0.52258807
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3fc526ca; // action129:  1.54024625
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h3fc51d2f; // action130:  1.53995311
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbfae5f44; // action131: -1.36228228
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h3fa6e0cc; // action132:  1.30373526
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3e23f410; // action133:  0.16011071
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3f2bfb5a; // action134:  0.67180407
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'hbe48f454; // action135: -0.19624454
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'hbfc6bc40; // action136: -1.55261993
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h3fe86958; // action137:  1.81571484
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h3ff19fe8; // action138:  1.88769245
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'h3fae6f02; // action139:  1.36276269
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'hbfa503cc; // action140: -1.28917837
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h3f98343f; // action141:  1.18909442
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3fec5650; // action142:  1.84638405
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'hbe76049c; // action143: -0.24025196
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'hbe36db6a; // action144: -0.17857137
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'hbee925e3; // action145: -0.45536718
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h3f9b75c7; // action146:  1.21453178
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbf87697d; // action147: -1.05790675
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3fdea85c; // action148:  1.73951292
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h3fcbcccf; // action149:  1.59218776
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'hbe32a3e9; // action150: -0.17445339
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbfd29869; // action151: -1.64527619
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3f8c651a; // action152:  1.09683537
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'hbf7ebaa1; // action153: -0.99503523
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h3ea0f912; // action154:  0.31440026
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'hbf9bbcac; // action155: -1.21669531
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbfda1dac; // action156: -1.70403051
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'h3fb180d2; // action157:  1.38674378
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'h3f9a31ba; // action158:  1.20464253
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h3f11a907; // action159:  0.56898540
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h3e73e443; // action160:  0.23817544
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'hbf84c0ce; // action161: -1.03713393
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'hbfe7f3d3; // action162: -1.81212842
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'hbfa54311; // action163: -1.29110920
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h3fd88d3d; // action164:  1.69181025
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'hbd116984; // action165: -0.03550102
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbead8748; // action166: -0.33892274
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbf8f6570; // action167: -1.12028313
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3f4647dd; // action168:  0.77453405
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbfd3ab7b; // action169: -1.65367067
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'h3f1f1604; // action170:  0.62142968
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'hbf6a8c68; // action171: -0.91620493
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3fd09f6d; // action172:  1.62986529
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'hbf210b54; // action173: -0.62907910
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'hbfa1e992; // action174: -1.26494050
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3f19c205; // action175:  0.60061675
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'hbf1bdb2a; // action176: -0.60881293
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'hbe19301e; // action177: -0.14959762
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbf03205a; // action178: -0.51221240
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h3f8e3e37; // action179:  1.11127365
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h3fb9b1a8; // action180:  1.45073414
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h3f442c57; // action181:  0.76630157
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbe1d9999; // action182: -0.15390624
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'hbfd33f7d; // action183: -1.65037501
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3fffb697; // action184:  1.99775970
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbf684101; // action185: -0.90724188
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'hbe7bf733; // action186: -0.24606018
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h3e9cd21c; // action187:  0.30629051
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'hbe83beb3; // action188: -0.25731429
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbf12a84b; // action189: -0.57288045
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h3fcd5813; // action190:  1.60425031
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h3edb4413; // action191:  0.42825374

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 16:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbe5eaf0c; // action0: -0.21746463
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3fcb1f18; // action1:  1.58688641
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3fed075a; // action2:  1.85178685
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'hbf471074; // action3: -0.77759480
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3f3bef75; // action4:  0.73412257
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h3fa2e8e5; // action5:  1.27273238
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'hbfdab018; // action6: -1.70849895
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h3f53d318; // action7:  0.82743979
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h3e28cc17; // action8:  0.16484104
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h3f4369d6; // action9:  0.76333368
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h3fc72b32; // action10:  1.55600572
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbd30eb0c; // action11: -0.04319291
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h3f67fa02; // action12:  0.90615857
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbfd147de; // action13: -1.63500571
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbf429390; // action14: -0.76006413
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3f2f3280; // action15:  0.68436432
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'hbf8cacc9; // action16: -1.09902298
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'hbfee588d; // action17: -1.86207736
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'hbe0394a4; // action18: -0.12849671
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'h3f0ecbb9; // action19:  0.55779606
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'hbf874ff6; // action20: -1.05712771
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbfb97252; // action21: -1.44880128
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h3f5b75d9; // action22:  0.85726696
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbfb61b2f; // action23: -1.42270458
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbf315ea7; // action24: -0.69285053
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3ff5fd27; // action25:  1.92178810
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h3fec1a5a; // action26:  1.84455419
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3fef1fdf; // action27:  1.86816013
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3f0021cc; // action28:  0.50051570
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbe3c76ae; // action29: -0.18404648
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'hbfb6454d; // action30: -1.42398989
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'h3f3530ce; // action31:  0.70777595
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbf95d601; // action32: -1.17059338
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3f0a7b5d; // action33:  0.54094487
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h3fbd0045; // action34:  1.47657073
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3f9c8ec1; // action35:  1.22310650
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3fadd879; // action36:  1.35816872
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h3ff61978; // action37:  1.92265224
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbf2528ad; // action38: -0.64515191
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'hbf9946b8; // action39: -1.19747066
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3ff84005; // action40:  1.93945372
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbecde079; // action41: -0.40210322
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'hbf9d2367; // action42: -1.22764289
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbf9e9476; // action43: -1.23890567
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3fc67c50; // action44:  1.55066872
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3f9dcd9d; // action45:  1.23283732
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h3f84324a; // action46:  1.03278470
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3fb02d2a; // action47:  1.37637830
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'hbedb0616; // action48: -0.42778081
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h3e213246; // action49:  0.15741834
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbff27e2a; // action50: -1.89447522
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbfe54e51; // action51: -1.79145253
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'h3f04efb9; // action52:  0.51928288
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h3fe023b5; // action53:  1.75108969
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'h3fa82512; // action54:  1.31363130
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'hbe3589fb; // action55: -0.17728417
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'h3fcb8706; // action56:  1.59005809
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbfe2594d; // action57: -1.76835024
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'hbffb2368; // action58: -1.96201801
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h3cc36ba5; // action59:  0.02385504
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbe740fdc; // action60: -0.23834175
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'hbf9f51d1; // action61: -1.24468434
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'h3f73f55f; // action62:  0.95296282
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3fd304c2; // action63:  1.64858270
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3fc849e2; // action64:  1.56475472
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3faf00b5; // action65:  1.36720908
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'hbfc870c7; // action66: -1.56594169
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbef8ccf6; // action67: -0.48593873
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3fa00c5a; // action68:  1.25037694
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3ea9959c; // action69:  0.33121955
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'hbeec674e; // action70: -0.46172565
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3fa742f0; // action71:  1.30673027
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3f09ceca; // action72:  0.53831160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3ff29eaa; // action73:  1.89546704
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3f396f0d; // action74:  0.72435075
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'hbed30103; // action75: -0.41211709
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'hbd27aec6; // action76: -0.04093816
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'h3fa208f2; // action77:  1.26589799
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h3f3627ea; // action78:  0.71154654
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h3ffb1384; // action79:  1.96153307
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'hbf95fa12; // action80: -1.17169404
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'hbf94222f; // action81: -1.15729320
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'hbfda06c3; // action82: -1.70333135
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'hbf718597; // action83: -0.94344467
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbfc06b88; // action84: -1.50328159
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbe094127; // action85: -0.13403760
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'hbfc2ecce; // action86: -1.52285171
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'hbf60cc66; // action87: -0.87811887
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbf72161d; // action88: -0.94564992
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h3efcc20c; // action89:  0.49366796
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3da185a8; // action90:  0.07886821
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3f3dfbec; // action91:  0.74212527
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h3e5eeca4; // action92:  0.21769959
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'hbfac7478; // action93: -1.34730434
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'hbff448c1; // action94: -1.90847027
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'h3f6e52c3; // action95:  0.93095034
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'h3fec12b5; // action96:  1.84432089
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'hbe0a111b; // action97: -0.13483088
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbebe25ee; // action98: -0.37138313
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3fa37000; // action99:  1.27685547
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'hbf8e63ab; // action100: -1.11241663
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h3eef6ab2; // action101:  0.46761090
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'hbf12e1e5; // action102: -0.57375938
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h3fd9b009; // action103:  1.70068467
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h3ff7736b; // action104:  1.93320978
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'h3fa9b1f7; // action105:  1.32574356
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3f95f4fe; // action106:  1.17153907
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbf896868; // action107: -1.07349873
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3f334731; // action108:  0.70030504
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'hbfc44beb; // action109: -1.53356683
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h3b6694ca; // action110:  0.00351839
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h3c47cd13; // action111:  0.01219489
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3f852bf2; // action112:  1.04040360
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h3fe0acb0; // action113:  1.75527000
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'hbfd13a9d; // action114: -1.63460124
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'hbeb7a684; // action115: -0.35869229
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3fc84fbc; // action116:  1.56493330
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3f45358e; // action117:  0.77034843
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3f29f6fb; // action118:  0.66392487
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3eec90d9; // action119:  0.46204260
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h3fe3b11a; // action120:  1.77884221
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3fd9de8d; // action121:  1.70210421
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'hbf207c0a; // action122: -0.62689269
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3e9509ed; // action123:  0.29109135
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'hbfda86ee; // action124: -1.70724273
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'hbfd3f25c; // action125: -1.65583372
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbed4266c; // action126: -0.41435564
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3fe38261; // action127:  1.77741635
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'h3f553feb; // action128:  0.83300656
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'hbf68e867; // action129: -0.90979618
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h3f468e04; // action130:  0.77560449
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h3ee66054; // action131:  0.44995368
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'h3fe10776; // action132:  1.75804019
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'hbf37b1cf; // action133: -0.71755689
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3f1b7841; // action134:  0.60730368
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h3ff151fb; // action135:  1.88531435
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h3fa512d0; // action136:  1.28963661
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h3e10330e; // action137:  0.14081976
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'hbf121531; // action138: -0.57063586
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'hbec49b78; // action139: -0.38399863
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'hbf3639c2; // action140: -0.71181881
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h3f4b2f08; // action141:  0.79368639
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3fd2e09e; // action142:  1.64747977
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h3f3b6997; // action143:  0.73207992
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'hbff92021; // action144: -1.94629300
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'hbf8063ae; // action145: -1.00304198
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h3f882da3; // action146:  1.06389272
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbfbaf8c2; // action147: -1.46071649
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3f2a238f; // action148:  0.66460508
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbfa48a3e; // action149: -1.28546882
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h3efb79f1; // action150:  0.49116471
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbfa0c056; // action151: -1.25586963
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'hbfbc6bd1; // action152: -1.47204030
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3f6b60fb; // action153:  0.91944855
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'hbe36b618; // action154: -0.17842901
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'hbdcdd488; // action155: -0.10050303
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'h3fcc3e27; // action156:  1.59564674
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbf2fcf3d; // action157: -0.68675596
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbfd34278; // action158: -1.65046597
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h3f8f8cda; // action159:  1.12148595
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbf920cfb; // action160: -1.14102113
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h3f5e9e97; // action161:  0.86960739
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h3f0c1aa7; // action162:  0.54728168
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h3fe53bf3; // action163:  1.79089200
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h3e3ec4a4; // action164:  0.18629700
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3f9efee3; // action165:  1.24215353
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbf52c28f; // action166: -0.82328123
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h3ff8ef12; // action167:  1.94479585
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3f07d485; // action168:  0.53058654
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h3f2c9c51; // action169:  0.67426020
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbe942f25; // action170: -0.28942218
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'hbc8df65d; // action171: -0.01732939
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'hbdb074ad; // action172: -0.08616004
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3f2a5092; // action173:  0.66529191
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3fad22e3; // action174:  1.35262716
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3ef79340; // action175:  0.48354530
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3fc35ce1; // action176:  1.52627194
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'hbf914a34; // action177: -1.13507700
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbf33d4fb; // action178: -0.70246857
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbf13b33a; // action179: -0.57695353
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'hbfb61429; // action180: -1.42249024
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h3f9b31b5; // action181:  1.21245444
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'h3fc8b6fa; // action182:  1.56808400
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'hbfc4f801; // action183: -1.53881848
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3fd02395; // action184:  1.62608588
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbe11d4fa; // action185: -0.14241400
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3fe135ae; // action186:  1.75945067
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'hbf449b56; // action187: -0.76799524
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h3ef1ddbb; // action188:  0.47239479
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbf6218f9; // action189: -0.88319355
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h3fbe5c92; // action190:  1.48720002
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h3fdf3ab1; // action191:  1.74397862

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 17:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'hbfaab176; // action0: -1.33354068
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3f44f7ce; // action1:  0.76940620
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'hbe431874; // action2: -0.19052297
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3ff30862; // action3:  1.89869332
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3fa24850; // action4:  1.26783180
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbf288400; // action5: -0.65826416
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3e97bdda; // action6:  0.29637033
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h3fdb7af8; // action7:  1.71469021
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h3fdfd83d; // action8:  1.74878657
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h3f95d33e; // action9:  1.17050910
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'h3fc5afd6; // action10:  1.54442859
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbf114cc7; // action11: -0.56757778
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'h3d7f45f6; // action12:  0.06232258
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbfc92589; // action13: -1.57145798
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbf6073e0; // action14: -0.87676811
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'hbf0e2d77; // action15: -0.55538124
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h3f867ebd; // action16:  1.05074275
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h3e9a7a2b; // action17:  0.30171332
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'hbfdfe735; // action18: -1.74924338
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbf6678be; // action19: -0.90027988
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'h3f83f8dd; // action20:  1.03103220
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbd65c036; // action21: -0.05609151
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'h3ee2b664; // action22:  0.44279778
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h3fd84b56; // action23:  1.68979907
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbff8979b; // action24: -1.94212663
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'hbfa8520c; // action25: -1.31500387
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'h3f7dec9b; // action26:  0.99189156
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'hbffd577d; // action27: -1.97923243
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3f767dd3; // action28:  0.96285743
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbe6ccd2c; // action29: -0.23125142
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3f7c6752; // action30:  0.98595154
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbed06094; // action31: -0.40698683
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h3f910157; // action32:  1.13285339
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'hbfb02de7; // action33: -1.37640083
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h3fb513ac; // action34:  1.41466284
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'hbfa37a9c; // action35: -1.27717924
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'hbfd59380; // action36: -1.66856384
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'hbfd1c199; // action37: -1.63872063
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h3fb7d323; // action38:  1.43613088
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h3e140513; // action39:  0.14455061
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3f8996de; // action40:  1.07491660
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h3fac8daf; // action41:  1.34807384
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3f58b7d3; // action42:  0.84655493
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbff78173; // action43: -1.93363798
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3f5cbaa6; // action44:  0.86222303
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'hbdab238e; // action45: -0.08356391
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h3e72078b; // action46:  0.23635690
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'h3f95a87f; // action47:  1.16920459
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'hbf02a5c5; // action48: -0.51034194
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h3f805f08; // action49:  1.00290012
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbfef28f0; // action50: -1.86843681
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h3f788f86; // action51:  0.97093999
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbfa930b7; // action52: -1.32179916
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'hbf341e65; // action53: -0.70358878
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'hbf108d75; // action54: -0.56465846
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h3fa0cc0b; // action55:  1.25622690
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'hbebcd606; // action56: -0.36882037
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbfd11cce; // action57: -1.63369155
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3e2d1f04; // action58:  0.16906363
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'hbe92ff2e; // action59: -0.28710312
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h3e740c85; // action60:  0.23832901
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'hbf845925; // action61: -1.03397048
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'hbfd0ebb5; // action62: -1.63219321
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3fb65d66; // action63:  1.42472529
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'h3ff0fcb8; // action64:  1.88271236
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'hbf83904e; // action65: -1.02784133
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h3fd145f3; // action66:  1.63494718
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbe9d497a; // action67: -0.30720121
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'hbee1fdfe; // action68: -0.44139093
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3fa9618e; // action69:  1.32328963
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'h3f833b13; // action70:  1.02524030
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3f769417; // action71:  0.96319717
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3ff01b1c; // action72:  1.87582731
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3df3f42e; // action73:  0.11911808
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3ffb9b56; // action74:  1.96567798
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3fc57674; // action75:  1.54267740
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h3fe12ae4; // action76:  1.75912142
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbf4712ea; // action77: -0.77763236
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h3f808e07; // action78:  1.00433433
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'hbe8a2030; // action79: -0.26977682
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'hbf37ac79; // action80: -0.71747547
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3fed857f; // action81:  1.85563648
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'hbf856da3; // action82: -1.04240835
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h3cd57919; // action83:  0.02605872
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'h3db33dbd; // action84:  0.08752010
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'h3d5babbd; // action85:  0.05363058
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h3efcfa03; // action86:  0.49409494
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3f9b8787; // action87:  1.21507347
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbf22495d; // action88: -0.63393193
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbfeb8a71; // action89: -1.84016240
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3f9243ab; // action90:  1.14269006
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'hbf00bac5; // action91: -0.50284988
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbfec4178; // action92: -1.84574795
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'hbf4b2a2b; // action93: -0.79361218
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'hbed691f5; // action94: -0.41908231
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'hbd520c6d; // action95: -0.05128138
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'hbefcc5d9; // action96: -0.49369696
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'hbe9266d5; // action97: -0.28594080
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'h3dbb846b; // action98:  0.09156116
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'h3e36278a; // action99:  0.17788520
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'hbfc7499a; // action100: -1.55693364
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h3fc6b88f; // action101:  1.55250728
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3f9ba674; // action102:  1.21601725
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h3fb1a382; // action103:  1.38780236
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'hbed2822b; // action104: -0.41114935
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbf0914a7; // action105: -0.53547138
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'hbf8f5ba8; // action106: -1.11998463
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbf1075e6; // action107: -0.56429899
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'hbef44dee; // action108: -0.47715706
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3eb096ca; // action109:  0.34490043
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h3fcad767; // action110:  1.58469856
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbe50e88a; // action111: -0.20401207
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'hbfeba4d7; // action112: -1.84096801
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h3f92aa45; // action113:  1.14582121
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'hbe5b3660; // action114: -0.21407461
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'hbfe76b42; // action115: -1.80796075
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3fa6691d; // action116:  1.30008280
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3f92b91a; // action117:  1.14627385
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'hbfca52b6; // action118: -1.58064914
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3f8a0589; // action119:  1.07829392
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h3ff69983; // action120:  1.92655981
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'hbec4ea50; // action121: -0.38460016
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'hbfeec0c6; // action122: -1.86525798
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'hbf2ea7bd; // action123: -0.68224698
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3ebd9928; // action124:  0.37030911
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'hbf33dd79; // action125: -0.70259815
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h3f68c718; // action126:  0.90928793
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3f168331; // action127:  0.58793932
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'hbf55162f; // action128: -0.83236974
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'hbf8ba796; // action129: -1.09105182
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'hbfed3123; // action130: -1.85306203
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h3d43488a; // action131:  0.04767660
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'hbe82f388; // action132: -0.25576425
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'hbd9c1b3b; // action133: -0.07622381
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3ffa63dd; // action134:  1.95617259
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'hbf96b44d; // action135: -1.17737734
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h3d2af059; // action136:  0.04173312
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h3f65dcf2; // action137:  0.89790261
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'hbf1fa190; // action138: -0.62355900
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'hbffbda35; // action139: -1.96759665
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h3f8c4446; // action140:  1.09583354
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'hbfbe5d38; // action141: -1.48721981
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3f7af2cc; // action142:  0.98026729
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'hbf451ca1; // action143: -0.76996809
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3fd530c4; // action144:  1.66555071
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'h3e98af37; // action145:  0.29821178
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'h3fb3a5eb; // action146:  1.40350091
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h3fe700ba; // action147:  1.80470967
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'hbeaabae7; // action148: -0.33345720
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbf01b8f9; // action149: -0.50672871
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h3f885e6f; // action150:  1.06538188
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h3fb16966; // action151:  1.38602901
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'hbfd1e6f1; // action152: -1.63986027
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'h3fd4fc24; // action153:  1.66394472
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'h3ffd37e2; // action154:  1.97826791
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'hbbe1bb71; // action155: -0.00688880
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbe51e53c; // action156: -0.20497602
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbfc1b383; // action157: -1.51329076
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbf439018; // action158: -0.76391745
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h3f95d6db; // action159:  1.17061937
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h3f1301e2; // action160:  0.57424748
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h3f91d29d; // action161:  1.13923991
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'hbfff0c68; // action162: -1.99256611
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'h3f64aad1; // action163:  0.89323145
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'h3f8eca24; // action164:  1.11554384
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3dcca885; // action165:  0.09993080
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h3f94e366; // action166:  1.16318965
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbd3e38a0; // action167: -0.04644072
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'hbf764e34; // action168: -0.96213078
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h3ffca9e5; // action169:  1.97393477
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbfeda97e; // action170: -1.85673499
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'hbf88628c; // action171: -1.06550741
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3fbc665a; // action172:  1.47187352
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'hbf52087c; // action173: -0.82044196
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'h3ff5c604; // action174:  1.92010546
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3f90b4b1; // action175:  1.13051426
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3f978a42; // action176:  1.18390679
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'hbedfca43; // action177: -0.43709001
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'h3f609cde; // action178:  0.87739360
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbee44588; // action179: -0.44584298
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h3f9b6096; // action180:  1.21388507
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h3fce155f; // action181:  1.61002719
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbfffe338; // action182: -1.99912167
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'hbe465599; // action183: -0.19368590
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'hbffde530; // action184: -1.98355675
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbe60242f; // action185: -0.21888803
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'h3e8855f0; // action186:  0.26628065
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'hbfadbca4; // action187: -1.35731936
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h3fdd53aa; // action188:  1.72911572
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'h3ec38412; // action189:  0.38186699
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'h3f8cdbc1; // action190:  1.10045636
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'h3f3c3545; // action191:  0.73518783

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 18:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h3e5c76a3; // action0:  0.21529631
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'hbf9b913d; // action1: -1.21536982
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'h3f291e51; // action2:  0.66061884
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'h3fc91ac3; // action3:  1.57112920
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'h3ca72db1; // action4:  0.02040753
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'h3fa7ed7f; // action5:  1.31193531
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3f8e8ecf; // action6:  1.11373317
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'h3f06cb73; // action7:  0.52654189
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h3ffc8a7c; // action8:  1.97297621
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'hbe3b3fc1; // action9: -0.18286039
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'hbfa4d24f; // action10: -1.28766811
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'hbf0caaaf; // action11: -0.54947942
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'hbfb75297; // action12: -1.43220794
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'hbff0c28b; // action13: -1.88093698
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'h3fdfeafc; // action14:  1.74935865
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'hbfd0ca44; // action15: -1.63117266
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'h3fb4da98; // action16:  1.41292095
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h3fa88db6; // action17:  1.31682467
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'h3faaefc9; // action18:  1.33544266
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbfaefed7; // action19: -1.36715209
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'hbfcbcd1a; // action20: -1.59219670
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'h3fa6c83d; // action21:  1.30298579
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'hbfcbb2fc; // action22: -1.59139967
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'hbf81d84e; // action23: -1.01441360
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbf359b91; // action24: -0.70940500
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'h3fd9027b; // action25:  1.69538820
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'hbfc3e036; // action26: -1.53027987
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'h3fe86aec; // action27:  1.81576300
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3f42ca79; // action28:  0.76090199
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbfbae6ee; // action29: -1.46017241
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3f7524ab; // action30:  0.95759076
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbeb68a63; // action31: -0.35652456
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'hbebf8de9; // action32: -0.37412956
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3fe1e1b0; // action33:  1.76469994
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'h3f47bd08; // action34:  0.78022814
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'hbfe585f6; // action35: -1.79315066
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'hbdd8eb81; // action36: -0.10591794
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'hbf84f624; // action37: -1.03876162
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'h3f8420c8; // action38:  1.03225040
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'hbfe5d70e; // action39: -1.79562545
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'hbfa7586a; // action40: -1.30738568
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'h3fc3d807; // action41:  1.53003013
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'h3f375919; // action42:  0.71620327
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'h3fca2c01; // action43:  1.57946789
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'h3f1ba5b5; // action44:  0.60799724
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'hbfd1a959; // action45: -1.63798058
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'hbe88288d; // action46: -0.26593438
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'hbee62e0c; // action47: -0.44957006
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'hbf8d79f3; // action48: -1.10528409
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h3fa8608b; // action49:  1.31544626
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbe7914fe; // action50: -0.24324414
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'hbf7dda9b; // action51: -0.99161690
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbfdc3d74; // action52: -1.72062540
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'hbf97123f; // action53: -1.18024433
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'hbe5347cf; // action54: -0.20632862
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'hbef42191; // action55: -0.47681859
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'hbfe16dc7; // action56: -1.76116264
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbf9551c4; // action57: -1.16655779
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3e7b431b; // action58:  0.24537317
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'hbf92e343; // action59: -1.14756048
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'hbdca6dfb; // action60: -0.09884258
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3fcabdcd; // action61:  1.58391726
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'hbfa483b7; // action62: -1.28526962
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'h3ffeb6e5; // action63:  1.98995650
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'hbfd6bd30; // action64: -1.67764854
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'hbdf9c64a; // action65: -0.12196024
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h3df426fe; // action66:  0.11921500
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'h3fb6a818; // action67:  1.42700481
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3f6a6bb1; // action68:  0.91570574
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'h3f24880a; // action69:  0.64270079
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'hbee42ea5; // action70: -0.44566837
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3f4a5c88; // action71:  0.79047441
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'h3e824a82; // action72:  0.25447470
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'hbf9f671d; // action73: -1.24533427
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'hbfe72392; // action74: -1.80577302
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3fdf7723; // action75:  1.74582326
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h3fab482e; // action76:  1.33814025
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbeea80db; // action77: -0.45801434
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'h3e8e95d6; // action78:  0.27848691
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h3f955661; // action79:  1.16669858
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3fc60999; // action80:  1.54716790
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'hbfc28092; // action81: -1.51954865
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'hbd4b1aee; // action82: -0.04958623
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h3ed85825; // action83:  0.42254749
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbfd68eb1; // action84: -1.67622960
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbee2c119; // action85: -0.44287947
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h3f90f64b; // action86:  1.13251626
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'h3fdc603a; // action87:  1.72168660
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbf6c134b; // action88: -0.92216939
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'hbfec2e5c; // action89: -1.84516478
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'hbf9b11a2; // action90: -1.21147561
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'hbffd3785; // action91: -1.97825682
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'hbdeaa30d; // action92: -0.11456881
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'hbf660f50; // action93: -0.89867115
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'h3f806544; // action94:  1.00309038
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'hbf0538fa; // action95: -0.52040064
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'hbf9c1f45; // action96: -1.21970427
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'hbf6322bd; // action97: -0.88724881
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbf76261a; // action98: -0.96151888
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'hbed65e44; // action99: -0.41868794
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h3fce2795; // action100:  1.61058295
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h3eacc185; // action101:  0.33741394
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'h3ded2541; // action102:  0.11579371
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'hbf89e2b8; // action103: -1.07723141
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'h3f2cc65c; // action104:  0.67490172
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbfe181b6; // action105: -1.76177096
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3ebc877a; // action106:  0.36822110
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'hbff04ca2; // action107: -1.87733865
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'hbefb852f; // action108: -0.49125049
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'hbff0c876; // action109: -1.88111758
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h3f8dcf03; // action110:  1.10788000
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'h3eabb0a1; // action111:  0.33533195
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'hbf54b2cc; // action112: -0.83085322
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'hbf29cc69; // action113: -0.66327530
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h3f3694d1; // action114:  0.71320826
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3e35da64; // action115:  0.17759091
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'hbec271df; // action116: -0.37977502
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'h3ef72ea3; // action117:  0.48277768
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'h3f2d4730; // action118:  0.67686749
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'hbf850e5d; // action119: -1.03950083
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h3c2b5a57; // action120:  0.01045855
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'h3f1a6659; // action121:  0.60312420
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'h3e9b3710; // action122:  0.30315447
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'h3f2a19d1; // action123:  0.66445643
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'h3fd25e3a; // action124:  1.64350057
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'hbfa91574; // action125: -1.32096720
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'hbf723b37; // action126: -0.94621605
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'hbeda0764; // action127: -0.42583764
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'hbe5c08f2; // action128: -0.21487787
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3fc5719d; // action129:  1.54252970
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h3f7311f9; // action130:  0.94949299
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'hbfe66266; // action131: -1.79987788
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'hbe8d2f4e; // action132: -0.27575153
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3f972190; // action133:  1.18071175
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'hbfa2e50a; // action134: -1.27261472
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h3fd37ab1; // action135:  1.65218174
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'hbfca0d56; // action136: -1.57853198
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h3f806531; // action137:  1.00308812
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'hbfcc019a; // action138: -1.59379888
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'hbfa4820d; // action139: -1.28521883
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'h3e4f4f12; // action140:  0.20245007
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'h3f2f417d; // action141:  0.68459302
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'h3fa01330; // action142:  1.25058556
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'h3fe2288f; // action143:  1.76686275
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3f73f743; // action144:  0.95299166
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'hbf072fbb; // action145: -0.52807206
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'hbfd7fa5d; // action146: -1.68732798
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'h3fdab6e0; // action147:  1.70870590
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3fc32497; // action148:  1.52455413
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'hbffb1036; // action149: -1.96143222
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h3f319106; // action150:  0.69361913
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'hbf269b0b; // action151: -0.65080327
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'h3f8368de; // action152:  1.02663779
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'hbfcc478e; // action153: -1.59593368
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'hbfd23c26; // action154: -1.64246058
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'h3f48fd90; // action155:  0.78511906
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbf8ec627; // action156: -1.11542213
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbe17167b; // action157: -0.14754669
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbeffc23e; // action158: -0.49952883
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'h3fcacfe4; // action159:  1.58446932
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'h3f99ce07; // action160:  1.20159996
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h3f533bd3; // action161:  0.82513160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'hbe8545e9; // action162: -0.26029900
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'hbf9a5d2a; // action163: -1.20596814
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbebb275a; // action164: -0.36553460
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3fa5b867; // action165:  1.29469001
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'hbfe6d4e3; // action166: -1.80337179
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'h3f159c30; // action167:  0.58441448
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'h3ff01b90; // action168:  1.87584114
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'h3f5368ca; // action169:  0.82581770
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbf129fa6; // action170: -0.57274854
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3fd16b67; // action171:  1.63609016
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3f69b5f3; // action172:  0.91293257
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3e55f6c2; // action173:  0.20894912
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'hbde8710d; // action174: -0.11349688
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3e3f0889; // action175:  0.18655600
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3fb2e8f3; // action176:  1.39773405
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'hbeb42098; // action177: -0.35181117
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbe91af3d; // action178: -0.28454009
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'hbef5909e; // action179: -0.47961897
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'h3fbcdbe6; // action180:  1.47546077
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'hbf362dbd; // action181: -0.71163541
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbf26a2ce; // action182: -0.65092170
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h3e869878; // action183:  0.26288199
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3ed898b6; // action184:  0.42304009
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbff122c2; // action185: -1.88387322
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'hbebb3c5b; // action186: -0.36569485
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h3fd9917f; // action187:  1.69975269
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h3fa51f78; // action188:  1.29002285
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbfb03713; // action189: -1.37668073
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'hbff5bc92; // action190: -1.91981721
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'hbfa46c80; // action191: -1.28456116

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
        // round 19:
            #24000 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd384; ram_i_data1 = 32'h3faca85e; // action0:  1.34888816
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd385; ram_i_data1 = 32'h3f6ab240; // action1:  0.91678238
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd386; ram_i_data1 = 32'hbfdf03f6; // action2: -1.74230838
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd387; ram_i_data1 = 32'hbf60334a; // action3: -0.87578261
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd388; ram_i_data1 = 32'hbfc928a0; // action4: -1.57155228
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd389; ram_i_data1 = 32'hbff5b416; // action5: -1.91955829
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd390; ram_i_data1 = 32'h3fa9ffd5; // action6:  1.32811987
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd391; ram_i_data1 = 32'hbf1d1c7d; // action7: -0.61371595
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd392; ram_i_data1 = 32'h3ffff352; // action8:  1.99961305
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd393; ram_i_data1 = 32'h3fbe688d; // action9:  1.48756564
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd394; ram_i_data1 = 32'hbf518ca1; // action10: -0.81855208
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd395; ram_i_data1 = 32'h3f2ada00; // action11:  0.66738892
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd396; ram_i_data1 = 32'hbff5524b; // action12: -1.91657388
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd397; ram_i_data1 = 32'h3fbf9dec; // action13:  1.49700689
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd398; ram_i_data1 = 32'hbff1fc38; // action14: -1.89050961
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd399; ram_i_data1 = 32'h3f9412a8; // action15:  1.15681934
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd400; ram_i_data1 = 32'hbf21e1a9; // action16: -0.63234955
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd401; ram_i_data1 = 32'h3fceeae8; // action17:  1.61654377
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd402; ram_i_data1 = 32'hbf00d725; // action18: -0.50328285
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd403; ram_i_data1 = 32'hbe8fe73d; // action19: -0.28106108
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd404; ram_i_data1 = 32'hbd845cdb; // action20: -0.06463023
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd405; ram_i_data1 = 32'hbf67f412; // action21: -0.90606797
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd406; ram_i_data1 = 32'hbff5baf1; // action22: -1.91976750
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd407; ram_i_data1 = 32'h3f586796; // action23:  0.84533060
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd408; ram_i_data1 = 32'hbfa15dc0; // action24: -1.26067352
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd409; ram_i_data1 = 32'hbfaab914; // action25: -1.33377314
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd410; ram_i_data1 = 32'hbf4a0559; // action26: -0.78914410
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd411; ram_i_data1 = 32'hbf653483; // action27: -0.89533252
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd412; ram_i_data1 = 32'h3ecf15c3; // action28:  0.40446290
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd413; ram_i_data1 = 32'hbf5fdc13; // action29: -0.87445182
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd414; ram_i_data1 = 32'h3fa5733f; // action30:  1.29257953
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd415; ram_i_data1 = 32'hbfab325b; // action31: -1.33747423
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd416; ram_i_data1 = 32'h3e895e95; // action32:  0.26829973
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd417; ram_i_data1 = 32'h3fe2f67a; // action33:  1.77314687
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd418; ram_i_data1 = 32'hbf364721; // action34: -0.71202284
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd419; ram_i_data1 = 32'h3e81405f; // action35:  0.25244424
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd420; ram_i_data1 = 32'h3fca9d22; // action36:  1.58292031
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd421; ram_i_data1 = 32'h3e29d803; // action37:  0.16586308
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd422; ram_i_data1 = 32'hbfd494a8; // action38: -1.66078663
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd423; ram_i_data1 = 32'h3fba4ccc; // action39:  1.45546865
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd424; ram_i_data1 = 32'h3b911af0; // action40:  0.00442826
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd425; ram_i_data1 = 32'hbffdeb3b; // action41: -1.98374116
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd426; ram_i_data1 = 32'hbf51d4f2; // action42: -0.81965554
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd427; ram_i_data1 = 32'hbe9ece61; // action43: -0.31016830
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd428; ram_i_data1 = 32'hbf4efb90; // action44: -0.80852604
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd429; ram_i_data1 = 32'h3f9ae599; // action45:  1.21013176
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd430; ram_i_data1 = 32'h3f4afc38; // action46:  0.79291105
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd431; ram_i_data1 = 32'hbf96baab; // action47: -1.17757165
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd432; ram_i_data1 = 32'h3ff8921d; // action48:  1.94195902
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd433; ram_i_data1 = 32'h3feb7aa5; // action49:  1.83968031
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd434; ram_i_data1 = 32'hbfa6d107; // action50: -1.30325401
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd435; ram_i_data1 = 32'h3e8dc848; // action51:  0.27691865
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd436; ram_i_data1 = 32'hbd8f147b; // action52: -0.06986328
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd437; ram_i_data1 = 32'h3f1de975; // action53:  0.61684352
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd438; ram_i_data1 = 32'hbe6ca632; // action54: -0.23110273
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd439; ram_i_data1 = 32'h3f024087; // action55:  0.50879711
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd440; ram_i_data1 = 32'hbfb9a030; // action56: -1.45020103
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd441; ram_i_data1 = 32'hbfa12950; // action57: -1.25907326
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd442; ram_i_data1 = 32'h3eef7302; // action58:  0.46767431
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd443; ram_i_data1 = 32'h3ffb3de6; // action59:  1.96282649
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd444; ram_i_data1 = 32'h3eb3de6e; // action60:  0.35130638
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd445; ram_i_data1 = 32'h3fc4b9d7; // action61:  1.53692138
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd446; ram_i_data1 = 32'hbfee8fa5; // action62: -1.86375868
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd447; ram_i_data1 = 32'hbe387822; // action63: -0.18014577
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd448; ram_i_data1 = 32'hbe7a3e6a; // action64: -0.24437872
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd449; ram_i_data1 = 32'h3fe31817; // action65:  1.77417266
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd450; ram_i_data1 = 32'h3fc863ed; // action66:  1.56554949
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd451; ram_i_data1 = 32'hbfbe180e; // action67: -1.48510909
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd452; ram_i_data1 = 32'h3f950cc1; // action68:  1.16445172
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd453; ram_i_data1 = 32'hbf3dc680; // action69: -0.74131012
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd454; ram_i_data1 = 32'hbf47d83e; // action70: -0.78064334
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd455; ram_i_data1 = 32'h3ef8a1c0; // action71:  0.48560905
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd456; ram_i_data1 = 32'hbfc0c528; // action72: -1.50601673
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd457; ram_i_data1 = 32'h3fd93573; // action73:  1.69694364
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd458; ram_i_data1 = 32'h3f794ac3; // action74:  0.97379702
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd459; ram_i_data1 = 32'h3dbe148e; // action75:  0.09281264
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd460; ram_i_data1 = 32'h3f0e668a; // action76:  0.55625212
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd461; ram_i_data1 = 32'hbce1f7b2; // action77: -0.02758393
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd462; ram_i_data1 = 32'hbf299840; // action78: -0.66247940
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd463; ram_i_data1 = 32'h3fc2d37a; // action79:  1.52207875
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd464; ram_i_data1 = 32'h3ff86a04; // action80:  1.94073534
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd465; ram_i_data1 = 32'h3d478463; // action81:  0.04871024
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd466; ram_i_data1 = 32'hbf77acdb; // action82: -0.96748132
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd467; ram_i_data1 = 32'h3fafade4; // action83:  1.37249422
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd468; ram_i_data1 = 32'hbf08b464; // action84: -0.53400254
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd469; ram_i_data1 = 32'hbf2f0e16; // action85: -0.68380868
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd470; ram_i_data1 = 32'h3ea67ce4; // action86:  0.32517159
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd471; ram_i_data1 = 32'hbf30fb42; // action87: -0.69133389
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd472; ram_i_data1 = 32'hbf424f7f; // action88: -0.75902551
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd473; ram_i_data1 = 32'h3ff917f9; // action89:  1.94604409
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd474; ram_i_data1 = 32'h3f3b6ddb; // action90:  0.73214501
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd475; ram_i_data1 = 32'h3f0931fc; // action91:  0.53591895
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd476; ram_i_data1 = 32'h3e6a385c; // action92:  0.22873062
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd477; ram_i_data1 = 32'h3fd72ab0; // action93:  1.68099022
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd478; ram_i_data1 = 32'hbfaab754; // action94: -1.33371973
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd479; ram_i_data1 = 32'hbf6e0695; // action95: -0.92978793
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd480; ram_i_data1 = 32'hbf2036bb; // action96: -0.62583512
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd481; ram_i_data1 = 32'h3fe24176; // action97:  1.76762271
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd482; ram_i_data1 = 32'hbe476be4; // action98: -0.19474751
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd483; ram_i_data1 = 32'hbfc7a3ac; // action99: -1.55968237
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd484; ram_i_data1 = 32'h3e3ac36f; // action100:  0.18238614
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd485; ram_i_data1 = 32'h3fc67863; // action101:  1.55054891
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd486; ram_i_data1 = 32'hbff70bca; // action102: -1.93004727
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd487; ram_i_data1 = 32'h3ff2a598; // action103:  1.89567852
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd488; ram_i_data1 = 32'hbee07e11; // action104: -0.43846181
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd489; ram_i_data1 = 32'hbf40e725; // action105: -0.75352699
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd490; ram_i_data1 = 32'h3fefe053; // action106:  1.87403333
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd491; ram_i_data1 = 32'h3fca87e6; // action107:  1.58227229
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd492; ram_i_data1 = 32'h3feb16a1; // action108:  1.83662808
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd493; ram_i_data1 = 32'h3fd3179a; // action109:  1.64915776
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd494; ram_i_data1 = 32'h3fb98b26; // action110:  1.44955897
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd495; ram_i_data1 = 32'hbfa79da4; // action111: -1.30949831
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd496; ram_i_data1 = 32'h3e8cddaa; // action112:  0.27512866
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd497; ram_i_data1 = 32'h3fb77b4a; // action113:  1.43344998
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd498; ram_i_data1 = 32'h3e487c2c; // action114:  0.19578618
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd499; ram_i_data1 = 32'h3fe3339c; // action115:  1.77501249
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd500; ram_i_data1 = 32'h3f8d7828; // action116:  1.10522938
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd501; ram_i_data1 = 32'hbf6bda4e; // action117: -0.92129982
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd502; ram_i_data1 = 32'hbfe22b38; // action118: -1.76694393
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd503; ram_i_data1 = 32'h3f16cc3f; // action119:  0.58905405
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd504; ram_i_data1 = 32'h3f4d70d5; // action120:  0.80250293
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd505; ram_i_data1 = 32'hbff69679; // action121: -1.92646706
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd506; ram_i_data1 = 32'hbf16e4a9; // action122: -0.58942658
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd507; ram_i_data1 = 32'hbff906b5; // action123: -1.94551718
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd508; ram_i_data1 = 32'hbfee85bb; // action124: -1.86345613
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd509; ram_i_data1 = 32'hbf0b51ba; // action125: -0.54421580
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd510; ram_i_data1 = 32'h3f63689d; // action126:  0.88831502
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd511; ram_i_data1 = 32'h3f23f9ec; // action127:  0.64053226
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd512; ram_i_data1 = 32'hbe1043c0; // action128: -0.14088345
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd513; ram_i_data1 = 32'h3f41fd1a; // action129:  0.75776827
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd514; ram_i_data1 = 32'h3e123000; // action130:  0.14276123
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd515; ram_i_data1 = 32'h3ec72083; // action131:  0.38891992
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd516; ram_i_data1 = 32'hbcfbfdc2; // action132: -0.03076065
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd517; ram_i_data1 = 32'h3f306559; // action133:  0.68904644
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd518; ram_i_data1 = 32'h3f8525bd; // action134:  1.04021418
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd519; ram_i_data1 = 32'h3fcd6ce9; // action135:  1.60488617
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd520; ram_i_data1 = 32'h3f75da42; // action136:  0.96036160
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd521; ram_i_data1 = 32'h3fbcae08; // action137:  1.47406101
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd522; ram_i_data1 = 32'h3f71e331; // action138:  0.94487292
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd523; ram_i_data1 = 32'hbf1aa690; // action139: -0.60410404
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd524; ram_i_data1 = 32'hbf9e9d1c; // action140: -1.23916960
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd525; ram_i_data1 = 32'hbfb8eb00; // action141: -1.44467163
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd526; ram_i_data1 = 32'hbfa7b43a; // action142: -1.31018758
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd527; ram_i_data1 = 32'hbffcf2a4; // action143: -1.97615480
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd528; ram_i_data1 = 32'h3fcd6232; // action144:  1.60455918
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd529; ram_i_data1 = 32'hbea75437; // action145: -0.32681438
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd530; ram_i_data1 = 32'hbfe4e2b8; // action146: -1.78816891
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd531; ram_i_data1 = 32'hbfcfbe0f; // action147: -1.62298763
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd532; ram_i_data1 = 32'h3fb8d8ec; // action148:  1.44411993
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd533; ram_i_data1 = 32'h3feeea16; // action149:  1.86651874
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd534; ram_i_data1 = 32'h3feacd6c; // action150:  1.83439398
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd535; ram_i_data1 = 32'h3e0375b4; // action151:  0.12837869
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd536; ram_i_data1 = 32'hbf88de80; // action152: -1.06929016
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd537; ram_i_data1 = 32'hbeb8d1b0; // action153: -0.36097479
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd538; ram_i_data1 = 32'hbfebf168; // action154: -1.84330463
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd539; ram_i_data1 = 32'hbf96fc46; // action155: -1.17957377
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd540; ram_i_data1 = 32'hbf38e1fc; // action156: -0.72219825
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd541; ram_i_data1 = 32'hbf6c1fea; // action157: -0.92236197
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd542; ram_i_data1 = 32'hbe98528c; // action158: -0.29750478
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd543; ram_i_data1 = 32'hbff71349; // action159: -1.93027604
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd544; ram_i_data1 = 32'hbf333498; // action160: -0.70002127
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd545; ram_i_data1 = 32'h3fefbec8; // action161:  1.87300968
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd546; ram_i_data1 = 32'h3e898abc; // action162:  0.26863658
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd547; ram_i_data1 = 32'hbfece29c; // action163: -1.85066557
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd548; ram_i_data1 = 32'hbf0ef962; // action164: -0.55849278
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd549; ram_i_data1 = 32'h3fa1e961; // action165:  1.26493466
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd550; ram_i_data1 = 32'h3f107342; // action166:  0.56425869
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd551; ram_i_data1 = 32'hbfd9a0c5; // action167: -1.70021880
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd552; ram_i_data1 = 32'hbfdf189b; // action168: -1.74293840
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd553; ram_i_data1 = 32'hbfc7a02f; // action169: -1.55957592
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd554; ram_i_data1 = 32'hbfe9b4bb; // action170: -1.82582796
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd555; ram_i_data1 = 32'h3eccd0a6; // action171:  0.40002936
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd556; ram_i_data1 = 32'h3f04680b; // action172:  0.51721257
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd557; ram_i_data1 = 32'h3fd8128c; // action173:  1.68806601
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd558; ram_i_data1 = 32'hbed11623; // action174: -0.40837201
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd559; ram_i_data1 = 32'h3fec8205; // action175:  1.84771788
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd560; ram_i_data1 = 32'h3e86c4c2; // action176:  0.26321989
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd561; ram_i_data1 = 32'hbf812f7c; // action177: -1.00926161
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd562; ram_i_data1 = 32'hbe418773; // action178: -0.18899326
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd563; ram_i_data1 = 32'h3fc6d1a4; // action179:  1.55327272
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd564; ram_i_data1 = 32'hbfa7a3ed; // action180: -1.30969012
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd565; ram_i_data1 = 32'h3fcb46dd; // action181:  1.58810008
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd566; ram_i_data1 = 32'hbeaf563a; // action182: -0.34245473
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd567; ram_i_data1 = 32'h3f735f38; // action183:  0.95067167
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd568; ram_i_data1 = 32'h3fc4c245; // action184:  1.53717864
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd569; ram_i_data1 = 32'hbf819fc5; // action185: -1.01268828
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd570; ram_i_data1 = 32'hbf56666e; // action186: -0.83750045
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd571; ram_i_data1 = 32'h3f7132a7; // action187:  0.94217914
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd572; ram_i_data1 = 32'h3fecc0ae; // action188:  1.84963012
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd573; ram_i_data1 = 32'hbf0cca0e; // action189: -0.54995811
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd574; ram_i_data1 = 32'hbfb18671; // action190: -1.38691533
            #10    ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd575; ram_i_data1 = 32'hbfbae76b; // action191: -1.46018732

            #10 ram_i_wr1 = 1'b0; ram_i_addr1 = 32'd576; ram_i_data1 = 32'd1; new_round = 1'b1; // start flag
            #10 ram_i_wr1 = 1'b1; ram_i_addr1 = 32'd0;   ram_i_data1 = 32'd0; new_round = 1'b0;
    end

    // record observations
        integer fpga_ans;
        localparam FPGA_ANS_WD_NUM = SW_ENV_NUM*(u_Pipeline.DST_ENV_WD_NUM-2) +
                                     SW_ENV_NUM*u_Pipeline.RWD_WL/DATA_WL +
                                     SW_ENV_NUM/DATA_WL;
        initial begin
            $display($clog2(1));
            fpga_ans = $fopen("/data0/FPGA_GYM/verilog/Pendulum/Pendulum.srcs/sim_1/new/fpga_ans.txt", "w");
            #640000 $fclose(fpga_ans);
        end
        always @(posedge new_round or negedge rstn) begin
            if (~rstn) begin
                cycle_cnt <= `ALL1(64);
            end else begin: write_fpga_ans
                reg [DATA_WL : 0] i;
                cycle_cnt <= cycle_cnt + 1;
                if (cycle_cnt[63] == 0) begin // there has been some result in BRAM
                    $fwrite(fpga_ans, "Iteration %d:\n", cycle_cnt);
                    for (i = `ZERO($clog2(SW_ENV_NUM)+1); i < FPGA_ANS_WD_NUM; i = i + 1) begin
                        $fwrite(fpga_ans, "%h%h%h%h ",
                                        u_My_RAM.Memory[u_Pipeline.OUT_INIT_ADDR+i][ 7: 0],
                                        u_My_RAM.Memory[u_Pipeline.OUT_INIT_ADDR+i][15: 8],
                                        u_My_RAM.Memory[u_Pipeline.OUT_INIT_ADDR+i][23:16],
                                        u_My_RAM.Memory[u_Pipeline.OUT_INIT_ADDR+i][31:24]);
                    end
                    $fwrite(fpga_ans, "\n\n");
                end
            end
        end

    // connect ports
        // Pipeline inputs
            assign uut_i_data = ram_o_data2;
        // BRAM inputs
            assign ram_i_wr2   = ~&uut_o_wea;
            assign ram_i_addr2 = uut_o_addr[ADDR_WL-1:2];
            assign ram_i_data2 = uut_o_data;

    Pipeline #(.DATA_WL(DATA_WL), .ADDR_WL(ADDR_WL), .WEA_WL(WEA_WL), .SW_ENV_NUM(SW_ENV_NUM)) u_Pipeline(
        .i_clk  ( clk  ),
        .i_rstn ( rstn ),
        .i_data ( uut_i_data[DATA_WL-1:0] ),
        .o_data ( uut_o_data[DATA_WL-1:0] ),
        .o_addr ( uut_o_addr[ADDR_WL-1:0] ),
        .o_en   ( uut_o_en ),
        .o_wea  ( uut_o_wea[WEA_WL-1:0] ),
        .o_rstb ( uut_o_rstb )
    );
    My_RAM #(.ADDR_WIDTH(RAM_ADDR_WL), .DATA_WIDTH(DATA_WL)) u_My_RAM(
        .i_clk   ( clk ),
        .i_rstn  ( rstn ),
        .i_wr1   ( ram_i_wr1 ),
        .i_addr1 ( ram_i_addr1[RAM_ADDR_WL-1:0] ),
        .i_data1 ( ram_i_data1[DATA_WL-1:0] ),
        .o_data1 ( ram_o_data1[DATA_WL-1:0] ),
        .i_wr2   ( ram_i_wr2 ),
        .i_addr2 ( ram_i_addr2[RAM_ADDR_WL-1:0] ),
        .i_data2 ( ram_i_data2[DATA_WL-1:0] ),
        .o_data2 ( ram_o_data2[DATA_WL-1:0] )
    );

endmodule
